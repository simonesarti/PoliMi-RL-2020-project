library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity project_tb is
end project_tb;

architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 100 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst	                : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		        : std_logic := '0';
signal   mem_o_data,mem_i_data	: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		        : std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);

signal RAM: ram_type := (0 => std_logic_vector(to_unsigned( 4 , 8)),
						1 => std_logic_vector(to_unsigned( 13 , 8)),
						2 => std_logic_vector(to_unsigned( 22 , 8)),
						3 => std_logic_vector(to_unsigned( 31 , 8)),
						4 => std_logic_vector(to_unsigned( 37 , 8)),
						5 => std_logic_vector(to_unsigned( 45 , 8)),
						6 => std_logic_vector(to_unsigned( 77 , 8)),
						7 => std_logic_vector(to_unsigned( 91 , 8)),
						8 => std_logic_vector(to_unsigned( 42 , 8)),
						others => (others =>'0'));

component project_reti_logiche is
port (
	i_clk         : in  std_logic;
	i_start       : in  std_logic;
	i_rst         : in  std_logic;
	i_data        : in  std_logic_vector(7 downto 0);
	o_address     : out std_logic_vector(15 downto 0);
	o_done        : out std_logic;
	o_en          : out std_logic;
	o_we          : out std_logic;
	o_data        : out std_logic_vector (7 downto 0)
	);
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
		i_clk      	=> tb_clk,
		i_start       => tb_start,
		i_rst      	=> tb_rst,
		i_data    	=> mem_o_data,
		o_address  	=> mem_address,
		o_done      	=> tb_done,
		o_en   	=> enable_wire,
		o_we 		=> mem_we,
		o_data    	=> mem_i_data
		);

p_CLK_GEN : process is
begin
	wait for c_CLOCK_PERIOD/2;
	tb_clk <= not tb_clk;
end process p_CLK_GEN;
MEM : process(tb_clk)
variable numero_test : integer := 0; --aggiunto per i test
begin
	if tb_clk'event and tb_clk = '1' then
		if enable_wire = '1' then
			if mem_we = '1' then
				RAM(conv_integer(mem_address))  <= mem_i_data;
				mem_o_data                      <= mem_i_data after 1 ns;
			else
				mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
			end if;
		end if;
		--modifico ram
		if(tb_rst='1') then

			if(numero_test = 0) then
				RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),1 => std_logic_vector(to_unsigned( 53, 8)),2 => std_logic_vector(to_unsigned( 75, 8)),3 => std_logic_vector(to_unsigned( 104, 8)),4 => std_logic_vector(to_unsigned( 113, 8)),5 => std_logic_vector(to_unsigned( 15, 8)),6 => std_logic_vector(to_unsigned( 124, 8)),7 => std_logic_vector(to_unsigned( 10, 8)),8 => std_logic_vector(to_unsigned( 32, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 1) then
				RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),1 => std_logic_vector(to_unsigned( 0, 8)),2 => std_logic_vector(to_unsigned( 105, 8)),3 => std_logic_vector(to_unsigned( 113, 8)),4 => std_logic_vector(to_unsigned( 86, 8)),5 => std_logic_vector(to_unsigned( 8, 8)),6 => std_logic_vector(to_unsigned( 95, 8)),7 => std_logic_vector(to_unsigned( 67, 8)),8 => std_logic_vector(to_unsigned( 54, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 2) then
				RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),1 => std_logic_vector(to_unsigned( 109, 8)),2 => std_logic_vector(to_unsigned( 78, 8)),3 => std_logic_vector(to_unsigned( 91, 8)),4 => std_logic_vector(to_unsigned( 8, 8)),5 => std_logic_vector(to_unsigned( 65, 8)),6 => std_logic_vector(to_unsigned( 17, 8)),7 => std_logic_vector(to_unsigned( 27, 8)),8 => std_logic_vector(to_unsigned( 75, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 3) then
				RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),1 => std_logic_vector(to_unsigned( 114, 8)),2 => std_logic_vector(to_unsigned( 46, 8)),3 => std_logic_vector(to_unsigned( 41, 8)),4 => std_logic_vector(to_unsigned( 1, 8)),5 => std_logic_vector(to_unsigned( 74, 8)),6 => std_logic_vector(to_unsigned( 119, 8)),7 => std_logic_vector(to_unsigned( 98, 8)),8 => std_logic_vector(to_unsigned( 101, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 4) then
				RAM <= (0 => std_logic_vector(to_unsigned( 90, 8)),1 => std_logic_vector(to_unsigned( 34, 8)),2 => std_logic_vector(to_unsigned( 7, 8)),3 => std_logic_vector(to_unsigned( 50, 8)),4 => std_logic_vector(to_unsigned( 113, 8)),5 => std_logic_vector(to_unsigned( 97, 8)),6 => std_logic_vector(to_unsigned( 17, 8)),7 => std_logic_vector(to_unsigned( 27, 8)),8 => std_logic_vector(to_unsigned( 118, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 5) then
				RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),1 => std_logic_vector(to_unsigned( 57, 8)),2 => std_logic_vector(to_unsigned( 24, 8)),3 => std_logic_vector(to_unsigned( 5, 8)),4 => std_logic_vector(to_unsigned( 36, 8)),5 => std_logic_vector(to_unsigned( 1, 8)),6 => std_logic_vector(to_unsigned( 90, 8)),7 => std_logic_vector(to_unsigned( 105, 8)),8 => std_logic_vector(to_unsigned( 35, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 6) then
				RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),1 => std_logic_vector(to_unsigned( 61, 8)),2 => std_logic_vector(to_unsigned( 78, 8)),3 => std_logic_vector(to_unsigned( 54, 8)),4 => std_logic_vector(to_unsigned( 48, 8)),5 => std_logic_vector(to_unsigned( 111, 8)),6 => std_logic_vector(to_unsigned( 101, 8)),7 => std_logic_vector(to_unsigned( 119, 8)),8 => std_logic_vector(to_unsigned( 56, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 7) then
				RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),1 => std_logic_vector(to_unsigned( 9, 8)),2 => std_logic_vector(to_unsigned( 13, 8)),3 => std_logic_vector(to_unsigned( 31, 8)),4 => std_logic_vector(to_unsigned( 24, 8)),5 => std_logic_vector(to_unsigned( 38, 8)),6 => std_logic_vector(to_unsigned( 4, 8)),7 => std_logic_vector(to_unsigned( 67, 8)),8 => std_logic_vector(to_unsigned( 100, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 8) then
				RAM <= (0 => std_logic_vector(to_unsigned( 91, 8)),1 => std_logic_vector(to_unsigned( 54, 8)),2 => std_logic_vector(to_unsigned( 9, 8)),3 => std_logic_vector(to_unsigned( 47, 8)),4 => std_logic_vector(to_unsigned( 17, 8)),5 => std_logic_vector(to_unsigned( 104, 8)),6 => std_logic_vector(to_unsigned( 35, 8)),7 => std_logic_vector(to_unsigned( 28, 8)),8 => std_logic_vector(to_unsigned( 52, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 9) then
				RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),1 => std_logic_vector(to_unsigned( 17, 8)),2 => std_logic_vector(to_unsigned( 6, 8)),3 => std_logic_vector(to_unsigned( 29, 8)),4 => std_logic_vector(to_unsigned( 112, 8)),5 => std_logic_vector(to_unsigned( 65, 8)),6 => std_logic_vector(to_unsigned( 102, 8)),7 => std_logic_vector(to_unsigned( 37, 8)),8 => std_logic_vector(to_unsigned( 4, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 10) then
				RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),1 => std_logic_vector(to_unsigned( 121, 8)),2 => std_logic_vector(to_unsigned( 46, 8)),3 => std_logic_vector(to_unsigned( 31, 8)),4 => std_logic_vector(to_unsigned( 22, 8)),5 => std_logic_vector(to_unsigned( 13, 8)),6 => std_logic_vector(to_unsigned( 37, 8)),7 => std_logic_vector(to_unsigned( 26, 8)),8 => std_logic_vector(to_unsigned( 100, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 11) then
				RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),1 => std_logic_vector(to_unsigned( 82, 8)),2 => std_logic_vector(to_unsigned( 9, 8)),3 => std_logic_vector(to_unsigned( 24, 8)),4 => std_logic_vector(to_unsigned( 28, 8)),5 => std_logic_vector(to_unsigned( 4, 8)),6 => std_logic_vector(to_unsigned( 65, 8)),7 => std_logic_vector(to_unsigned( 53, 8)),8 => std_logic_vector(to_unsigned( 79, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 12) then
				RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),1 => std_logic_vector(to_unsigned( 26, 8)),2 => std_logic_vector(to_unsigned( 60, 8)),3 => std_logic_vector(to_unsigned( 72, 8)),4 => std_logic_vector(to_unsigned( 33, 8)),5 => std_logic_vector(to_unsigned( 113, 8)),6 => std_logic_vector(to_unsigned( 97, 8)),7 => std_logic_vector(to_unsigned( 3, 8)),8 => std_logic_vector(to_unsigned( 47, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 13) then
				RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),1 => std_logic_vector(to_unsigned( 11, 8)),2 => std_logic_vector(to_unsigned( 33, 8)),3 => std_logic_vector(to_unsigned( 88, 8)),4 => std_logic_vector(to_unsigned( 83, 8)),5 => std_logic_vector(to_unsigned( 97, 8)),6 => std_logic_vector(to_unsigned( 66, 8)),7 => std_logic_vector(to_unsigned( 73, 8)),8 => std_logic_vector(to_unsigned( 76, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 14) then
				RAM <= (0 => std_logic_vector(to_unsigned( 71, 8)),1 => std_logic_vector(to_unsigned( 48, 8)),2 => std_logic_vector(to_unsigned( 24, 8)),3 => std_logic_vector(to_unsigned( 31, 8)),4 => std_logic_vector(to_unsigned( 67, 8)),5 => std_logic_vector(to_unsigned( 93, 8)),6 => std_logic_vector(to_unsigned( 1, 8)),7 => std_logic_vector(to_unsigned( 76, 8)),8 => std_logic_vector(to_unsigned( 62, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 15) then
				RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),1 => std_logic_vector(to_unsigned( 77, 8)),2 => std_logic_vector(to_unsigned( 110, 8)),3 => std_logic_vector(to_unsigned( 106, 8)),4 => std_logic_vector(to_unsigned( 70, 8)),5 => std_logic_vector(to_unsigned( 18, 8)),6 => std_logic_vector(to_unsigned( 83, 8)),7 => std_logic_vector(to_unsigned( 38, 8)),8 => std_logic_vector(to_unsigned( 93, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 16) then
				RAM <= (0 => std_logic_vector(to_unsigned( 62, 8)),1 => std_logic_vector(to_unsigned( 41, 8)),2 => std_logic_vector(to_unsigned( 120, 8)),3 => std_logic_vector(to_unsigned( 96, 8)),4 => std_logic_vector(to_unsigned( 36, 8)),5 => std_logic_vector(to_unsigned( 70, 8)),6 => std_logic_vector(to_unsigned( 111, 8)),7 => std_logic_vector(to_unsigned( 57, 8)),8 => std_logic_vector(to_unsigned( 26, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 17) then
				RAM <= (0 => std_logic_vector(to_unsigned( 8, 8)),1 => std_logic_vector(to_unsigned( 3, 8)),2 => std_logic_vector(to_unsigned( 76, 8)),3 => std_logic_vector(to_unsigned( 122, 8)),4 => std_logic_vector(to_unsigned( 62, 8)),5 => std_logic_vector(to_unsigned( 87, 8)),6 => std_logic_vector(to_unsigned( 24, 8)),7 => std_logic_vector(to_unsigned( 41, 8)),8 => std_logic_vector(to_unsigned( 76, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 18) then
				RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),1 => std_logic_vector(to_unsigned( 48, 8)),2 => std_logic_vector(to_unsigned( 9, 8)),3 => std_logic_vector(to_unsigned( 68, 8)),4 => std_logic_vector(to_unsigned( 38, 8)),5 => std_logic_vector(to_unsigned( 123, 8)),6 => std_logic_vector(to_unsigned( 75, 8)),7 => std_logic_vector(to_unsigned( 80, 8)),8 => std_logic_vector(to_unsigned( 68, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 19) then
				RAM <= (0 => std_logic_vector(to_unsigned( 5, 8)),1 => std_logic_vector(to_unsigned( 20, 8)),2 => std_logic_vector(to_unsigned( 69, 8)),3 => std_logic_vector(to_unsigned( 96, 8)),4 => std_logic_vector(to_unsigned( 47, 8)),5 => std_logic_vector(to_unsigned( 84, 8)),6 => std_logic_vector(to_unsigned( 43, 8)),7 => std_logic_vector(to_unsigned( 36, 8)),8 => std_logic_vector(to_unsigned( 25, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 20) then
				RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),1 => std_logic_vector(to_unsigned( 45, 8)),2 => std_logic_vector(to_unsigned( 85, 8)),3 => std_logic_vector(to_unsigned( 114, 8)),4 => std_logic_vector(to_unsigned( 74, 8)),5 => std_logic_vector(to_unsigned( 102, 8)),6 => std_logic_vector(to_unsigned( 106, 8)),7 => std_logic_vector(to_unsigned( 60, 8)),8 => std_logic_vector(to_unsigned( 107, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 21) then
				RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),1 => std_logic_vector(to_unsigned( 115, 8)),2 => std_logic_vector(to_unsigned( 124, 8)),3 => std_logic_vector(to_unsigned( 65, 8)),4 => std_logic_vector(to_unsigned( 89, 8)),5 => std_logic_vector(to_unsigned( 59, 8)),6 => std_logic_vector(to_unsigned( 39, 8)),7 => std_logic_vector(to_unsigned( 44, 8)),8 => std_logic_vector(to_unsigned( 110, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 22) then
				RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),1 => std_logic_vector(to_unsigned( 32, 8)),2 => std_logic_vector(to_unsigned( 106, 8)),3 => std_logic_vector(to_unsigned( 77, 8)),4 => std_logic_vector(to_unsigned( 40, 8)),5 => std_logic_vector(to_unsigned( 99, 8)),6 => std_logic_vector(to_unsigned( 24, 8)),7 => std_logic_vector(to_unsigned( 28, 8)),8 => std_logic_vector(to_unsigned( 84, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 23) then
				RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),1 => std_logic_vector(to_unsigned( 6, 8)),2 => std_logic_vector(to_unsigned( 93, 8)),3 => std_logic_vector(to_unsigned( 119, 8)),4 => std_logic_vector(to_unsigned( 72, 8)),5 => std_logic_vector(to_unsigned( 50, 8)),6 => std_logic_vector(to_unsigned( 10, 8)),7 => std_logic_vector(to_unsigned( 124, 8)),8 => std_logic_vector(to_unsigned( 62, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 24) then
				RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),1 => std_logic_vector(to_unsigned( 37, 8)),2 => std_logic_vector(to_unsigned( 124, 8)),3 => std_logic_vector(to_unsigned( 101, 8)),4 => std_logic_vector(to_unsigned( 96, 8)),5 => std_logic_vector(to_unsigned( 91, 8)),6 => std_logic_vector(to_unsigned( 33, 8)),7 => std_logic_vector(to_unsigned( 8, 8)),8 => std_logic_vector(to_unsigned( 115, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 25) then
				RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),1 => std_logic_vector(to_unsigned( 1, 8)),2 => std_logic_vector(to_unsigned( 110, 8)),3 => std_logic_vector(to_unsigned( 101, 8)),4 => std_logic_vector(to_unsigned( 52, 8)),5 => std_logic_vector(to_unsigned( 58, 8)),6 => std_logic_vector(to_unsigned( 86, 8)),7 => std_logic_vector(to_unsigned( 19, 8)),8 => std_logic_vector(to_unsigned( 34, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 26) then
				RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),1 => std_logic_vector(to_unsigned( 31, 8)),2 => std_logic_vector(to_unsigned( 89, 8)),3 => std_logic_vector(to_unsigned( 116, 8)),4 => std_logic_vector(to_unsigned( 122, 8)),5 => std_logic_vector(to_unsigned( 51, 8)),6 => std_logic_vector(to_unsigned( 16, 8)),7 => std_logic_vector(to_unsigned( 45, 8)),8 => std_logic_vector(to_unsigned( 122, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 27) then
				RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),1 => std_logic_vector(to_unsigned( 98, 8)),2 => std_logic_vector(to_unsigned( 121, 8)),3 => std_logic_vector(to_unsigned( 89, 8)),4 => std_logic_vector(to_unsigned( 93, 8)),5 => std_logic_vector(to_unsigned( 63, 8)),6 => std_logic_vector(to_unsigned( 23, 8)),7 => std_logic_vector(to_unsigned( 70, 8)),8 => std_logic_vector(to_unsigned( 14, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 28) then
				RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),1 => std_logic_vector(to_unsigned( 122, 8)),2 => std_logic_vector(to_unsigned( 2, 8)),3 => std_logic_vector(to_unsigned( 9, 8)),4 => std_logic_vector(to_unsigned( 20, 8)),5 => std_logic_vector(to_unsigned( 76, 8)),6 => std_logic_vector(to_unsigned( 16, 8)),7 => std_logic_vector(to_unsigned( 103, 8)),8 => std_logic_vector(to_unsigned( 25, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 29) then
				RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),1 => std_logic_vector(to_unsigned( 113, 8)),2 => std_logic_vector(to_unsigned( 61, 8)),3 => std_logic_vector(to_unsigned( 82, 8)),4 => std_logic_vector(to_unsigned( 39, 8)),5 => std_logic_vector(to_unsigned( 92, 8)),6 => std_logic_vector(to_unsigned( 124, 8)),7 => std_logic_vector(to_unsigned( 26, 8)),8 => std_logic_vector(to_unsigned( 29, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 30) then
				RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),1 => std_logic_vector(to_unsigned( 58, 8)),2 => std_logic_vector(to_unsigned( 62, 8)),3 => std_logic_vector(to_unsigned( 54, 8)),4 => std_logic_vector(to_unsigned( 72, 8)),5 => std_logic_vector(to_unsigned( 82, 8)),6 => std_logic_vector(to_unsigned( 107, 8)),7 => std_logic_vector(to_unsigned( 86, 8)),8 => std_logic_vector(to_unsigned( 102, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 31) then
				RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),1 => std_logic_vector(to_unsigned( 48, 8)),2 => std_logic_vector(to_unsigned( 69, 8)),3 => std_logic_vector(to_unsigned( 29, 8)),4 => std_logic_vector(to_unsigned( 105, 8)),5 => std_logic_vector(to_unsigned( 55, 8)),6 => std_logic_vector(to_unsigned( 121, 8)),7 => std_logic_vector(to_unsigned( 41, 8)),8 => std_logic_vector(to_unsigned( 64, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 32) then
				RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),1 => std_logic_vector(to_unsigned( 6, 8)),2 => std_logic_vector(to_unsigned( 17, 8)),3 => std_logic_vector(to_unsigned( 37, 8)),4 => std_logic_vector(to_unsigned( 68, 8)),5 => std_logic_vector(to_unsigned( 2, 8)),6 => std_logic_vector(to_unsigned( 98, 8)),7 => std_logic_vector(to_unsigned( 32, 8)),8 => std_logic_vector(to_unsigned( 53, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 33) then
				RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),1 => std_logic_vector(to_unsigned( 101, 8)),2 => std_logic_vector(to_unsigned( 118, 8)),3 => std_logic_vector(to_unsigned( 94, 8)),4 => std_logic_vector(to_unsigned( 4, 8)),5 => std_logic_vector(to_unsigned( 80, 8)),6 => std_logic_vector(to_unsigned( 73, 8)),7 => std_logic_vector(to_unsigned( 84, 8)),8 => std_logic_vector(to_unsigned( 89, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 34) then
				RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),1 => std_logic_vector(to_unsigned( 32, 8)),2 => std_logic_vector(to_unsigned( 22, 8)),3 => std_logic_vector(to_unsigned( 77, 8)),4 => std_logic_vector(to_unsigned( 27, 8)),5 => std_logic_vector(to_unsigned( 81, 8)),6 => std_logic_vector(to_unsigned( 48, 8)),7 => std_logic_vector(to_unsigned( 99, 8)),8 => std_logic_vector(to_unsigned( 112, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 35) then
				RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),1 => std_logic_vector(to_unsigned( 19, 8)),2 => std_logic_vector(to_unsigned( 36, 8)),3 => std_logic_vector(to_unsigned( 85, 8)),4 => std_logic_vector(to_unsigned( 108, 8)),5 => std_logic_vector(to_unsigned( 14, 8)),6 => std_logic_vector(to_unsigned( 50, 8)),7 => std_logic_vector(to_unsigned( 55, 8)),8 => std_logic_vector(to_unsigned( 100, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 36) then
				RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),1 => std_logic_vector(to_unsigned( 63, 8)),2 => std_logic_vector(to_unsigned( 7, 8)),3 => std_logic_vector(to_unsigned( 0, 8)),4 => std_logic_vector(to_unsigned( 124, 8)),5 => std_logic_vector(to_unsigned( 77, 8)),6 => std_logic_vector(to_unsigned( 94, 8)),7 => std_logic_vector(to_unsigned( 68, 8)),8 => std_logic_vector(to_unsigned( 67, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 37) then
				RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),1 => std_logic_vector(to_unsigned( 14, 8)),2 => std_logic_vector(to_unsigned( 37, 8)),3 => std_logic_vector(to_unsigned( 27, 8)),4 => std_logic_vector(to_unsigned( 33, 8)),5 => std_logic_vector(to_unsigned( 21, 8)),6 => std_logic_vector(to_unsigned( 41, 8)),7 => std_logic_vector(to_unsigned( 70, 8)),8 => std_logic_vector(to_unsigned( 106, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 38) then
				RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),1 => std_logic_vector(to_unsigned( 110, 8)),2 => std_logic_vector(to_unsigned( 69, 8)),3 => std_logic_vector(to_unsigned( 9, 8)),4 => std_logic_vector(to_unsigned( 47, 8)),5 => std_logic_vector(to_unsigned( 85, 8)),6 => std_logic_vector(to_unsigned( 19, 8)),7 => std_logic_vector(to_unsigned( 65, 8)),8 => std_logic_vector(to_unsigned( 65, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 39) then
				RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),1 => std_logic_vector(to_unsigned( 7, 8)),2 => std_logic_vector(to_unsigned( 95, 8)),3 => std_logic_vector(to_unsigned( 51, 8)),4 => std_logic_vector(to_unsigned( 71, 8)),5 => std_logic_vector(to_unsigned( 33, 8)),6 => std_logic_vector(to_unsigned( 56, 8)),7 => std_logic_vector(to_unsigned( 1, 8)),8 => std_logic_vector(to_unsigned( 107, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 40) then
				RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),1 => std_logic_vector(to_unsigned( 96, 8)),2 => std_logic_vector(to_unsigned( 52, 8)),3 => std_logic_vector(to_unsigned( 69, 8)),4 => std_logic_vector(to_unsigned( 59, 8)),5 => std_logic_vector(to_unsigned( 116, 8)),6 => std_logic_vector(to_unsigned( 104, 8)),7 => std_logic_vector(to_unsigned( 29, 8)),8 => std_logic_vector(to_unsigned( 46, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 41) then
				RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),1 => std_logic_vector(to_unsigned( 66, 8)),2 => std_logic_vector(to_unsigned( 105, 8)),3 => std_logic_vector(to_unsigned( 80, 8)),4 => std_logic_vector(to_unsigned( 72, 8)),5 => std_logic_vector(to_unsigned( 51, 8)),6 => std_logic_vector(to_unsigned( 36, 8)),7 => std_logic_vector(to_unsigned( 28, 8)),8 => std_logic_vector(to_unsigned( 35, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 42) then
				RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),1 => std_logic_vector(to_unsigned( 64, 8)),2 => std_logic_vector(to_unsigned( 120, 8)),3 => std_logic_vector(to_unsigned( 28, 8)),4 => std_logic_vector(to_unsigned( 94, 8)),5 => std_logic_vector(to_unsigned( 15, 8)),6 => std_logic_vector(to_unsigned( 49, 8)),7 => std_logic_vector(to_unsigned( 77, 8)),8 => std_logic_vector(to_unsigned( 56, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 43) then
				RAM <= (0 => std_logic_vector(to_unsigned( 70, 8)),1 => std_logic_vector(to_unsigned( 28, 8)),2 => std_logic_vector(to_unsigned( 116, 8)),3 => std_logic_vector(to_unsigned( 21, 8)),4 => std_logic_vector(to_unsigned( 86, 8)),5 => std_logic_vector(to_unsigned( 13, 8)),6 => std_logic_vector(to_unsigned( 64, 8)),7 => std_logic_vector(to_unsigned( 33, 8)),8 => std_logic_vector(to_unsigned( 41, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 44) then
				RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),1 => std_logic_vector(to_unsigned( 92, 8)),2 => std_logic_vector(to_unsigned( 108, 8)),3 => std_logic_vector(to_unsigned( 15, 8)),4 => std_logic_vector(to_unsigned( 66, 8)),5 => std_logic_vector(to_unsigned( 73, 8)),6 => std_logic_vector(to_unsigned( 102, 8)),7 => std_logic_vector(to_unsigned( 33, 8)),8 => std_logic_vector(to_unsigned( 23, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 45) then
				RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),1 => std_logic_vector(to_unsigned( 25, 8)),2 => std_logic_vector(to_unsigned( 16, 8)),3 => std_logic_vector(to_unsigned( 108, 8)),4 => std_logic_vector(to_unsigned( 113, 8)),5 => std_logic_vector(to_unsigned( 0, 8)),6 => std_logic_vector(to_unsigned( 102, 8)),7 => std_logic_vector(to_unsigned( 61, 8)),8 => std_logic_vector(to_unsigned( 62, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 46) then
				RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),1 => std_logic_vector(to_unsigned( 124, 8)),2 => std_logic_vector(to_unsigned( 58, 8)),3 => std_logic_vector(to_unsigned( 95, 8)),4 => std_logic_vector(to_unsigned( 29, 8)),5 => std_logic_vector(to_unsigned( 66, 8)),6 => std_logic_vector(to_unsigned( 12, 8)),7 => std_logic_vector(to_unsigned( 54, 8)),8 => std_logic_vector(to_unsigned( 126, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 47) then
				RAM <= (0 => std_logic_vector(to_unsigned( 4, 8)),1 => std_logic_vector(to_unsigned( 72, 8)),2 => std_logic_vector(to_unsigned( 53, 8)),3 => std_logic_vector(to_unsigned( 76, 8)),4 => std_logic_vector(to_unsigned( 110, 8)),5 => std_logic_vector(to_unsigned( 39, 8)),6 => std_logic_vector(to_unsigned( 49, 8)),7 => std_logic_vector(to_unsigned( 91, 8)),8 => std_logic_vector(to_unsigned( 55, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 48) then
				RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),1 => std_logic_vector(to_unsigned( 96, 8)),2 => std_logic_vector(to_unsigned( 74, 8)),3 => std_logic_vector(to_unsigned( 57, 8)),4 => std_logic_vector(to_unsigned( 101, 8)),5 => std_logic_vector(to_unsigned( 19, 8)),6 => std_logic_vector(to_unsigned( 112, 8)),7 => std_logic_vector(to_unsigned( 124, 8)),8 => std_logic_vector(to_unsigned( 27, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 49) then
				RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),1 => std_logic_vector(to_unsigned( 0, 8)),2 => std_logic_vector(to_unsigned( 36, 8)),3 => std_logic_vector(to_unsigned( 112, 8)),4 => std_logic_vector(to_unsigned( 87, 8)),5 => std_logic_vector(to_unsigned( 102, 8)),6 => std_logic_vector(to_unsigned( 92, 8)),7 => std_logic_vector(to_unsigned( 124, 8)),8 => std_logic_vector(to_unsigned( 116, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 50) then
				RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),1 => std_logic_vector(to_unsigned( 16, 8)),2 => std_logic_vector(to_unsigned( 79, 8)),3 => std_logic_vector(to_unsigned( 69, 8)),4 => std_logic_vector(to_unsigned( 118, 8)),5 => std_logic_vector(to_unsigned( 8, 8)),6 => std_logic_vector(to_unsigned( 53, 8)),7 => std_logic_vector(to_unsigned( 94, 8)),8 => std_logic_vector(to_unsigned( 81, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 51) then
				RAM <= (0 => std_logic_vector(to_unsigned( 47, 8)),1 => std_logic_vector(to_unsigned( 57, 8)),2 => std_logic_vector(to_unsigned( 35, 8)),3 => std_logic_vector(to_unsigned( 40, 8)),4 => std_logic_vector(to_unsigned( 118, 8)),5 => std_logic_vector(to_unsigned( 108, 8)),6 => std_logic_vector(to_unsigned( 65, 8)),7 => std_logic_vector(to_unsigned( 80, 8)),8 => std_logic_vector(to_unsigned( 72, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 52) then
				RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),1 => std_logic_vector(to_unsigned( 114, 8)),2 => std_logic_vector(to_unsigned( 49, 8)),3 => std_logic_vector(to_unsigned( 78, 8)),4 => std_logic_vector(to_unsigned( 4, 8)),5 => std_logic_vector(to_unsigned( 73, 8)),6 => std_logic_vector(to_unsigned( 92, 8)),7 => std_logic_vector(to_unsigned( 20, 8)),8 => std_logic_vector(to_unsigned( 79, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 53) then
				RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),1 => std_logic_vector(to_unsigned( 116, 8)),2 => std_logic_vector(to_unsigned( 85, 8)),3 => std_logic_vector(to_unsigned( 67, 8)),4 => std_logic_vector(to_unsigned( 46, 8)),5 => std_logic_vector(to_unsigned( 38, 8)),6 => std_logic_vector(to_unsigned( 23, 8)),7 => std_logic_vector(to_unsigned( 111, 8)),8 => std_logic_vector(to_unsigned( 113, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 54) then
				RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),1 => std_logic_vector(to_unsigned( 65, 8)),2 => std_logic_vector(to_unsigned( 27, 8)),3 => std_logic_vector(to_unsigned( 45, 8)),4 => std_logic_vector(to_unsigned( 40, 8)),5 => std_logic_vector(to_unsigned( 17, 8)),6 => std_logic_vector(to_unsigned( 84, 8)),7 => std_logic_vector(to_unsigned( 23, 8)),8 => std_logic_vector(to_unsigned( 84, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 55) then
				RAM <= (0 => std_logic_vector(to_unsigned( 70, 8)),1 => std_logic_vector(to_unsigned( 82, 8)),2 => std_logic_vector(to_unsigned( 64, 8)),3 => std_logic_vector(to_unsigned( 26, 8)),4 => std_logic_vector(to_unsigned( 6, 8)),5 => std_logic_vector(to_unsigned( 117, 8)),6 => std_logic_vector(to_unsigned( 113, 8)),7 => std_logic_vector(to_unsigned( 49, 8)),8 => std_logic_vector(to_unsigned( 59, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 56) then
				RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),1 => std_logic_vector(to_unsigned( 32, 8)),2 => std_logic_vector(to_unsigned( 24, 8)),3 => std_logic_vector(to_unsigned( 88, 8)),4 => std_logic_vector(to_unsigned( 28, 8)),5 => std_logic_vector(to_unsigned( 4, 8)),6 => std_logic_vector(to_unsigned( 43, 8)),7 => std_logic_vector(to_unsigned( 14, 8)),8 => std_logic_vector(to_unsigned( 99, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 57) then
				RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),1 => std_logic_vector(to_unsigned( 4, 8)),2 => std_logic_vector(to_unsigned( 110, 8)),3 => std_logic_vector(to_unsigned( 38, 8)),4 => std_logic_vector(to_unsigned( 122, 8)),5 => std_logic_vector(to_unsigned( 12, 8)),6 => std_logic_vector(to_unsigned( 95, 8)),7 => std_logic_vector(to_unsigned( 61, 8)),8 => std_logic_vector(to_unsigned( 94, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 58) then
				RAM <= (0 => std_logic_vector(to_unsigned( 4, 8)),1 => std_logic_vector(to_unsigned( 88, 8)),2 => std_logic_vector(to_unsigned( 105, 8)),3 => std_logic_vector(to_unsigned( 56, 8)),4 => std_logic_vector(to_unsigned( 81, 8)),5 => std_logic_vector(to_unsigned( 34, 8)),6 => std_logic_vector(to_unsigned( 97, 8)),7 => std_logic_vector(to_unsigned( 110, 8)),8 => std_logic_vector(to_unsigned( 124, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 59) then
				RAM <= (0 => std_logic_vector(to_unsigned( 46, 8)),1 => std_logic_vector(to_unsigned( 88, 8)),2 => std_logic_vector(to_unsigned( 101, 8)),3 => std_logic_vector(to_unsigned( 27, 8)),4 => std_logic_vector(to_unsigned( 83, 8)),5 => std_logic_vector(to_unsigned( 37, 8)),6 => std_logic_vector(to_unsigned( 55, 8)),7 => std_logic_vector(to_unsigned( 15, 8)),8 => std_logic_vector(to_unsigned( 31, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 60) then
				RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),1 => std_logic_vector(to_unsigned( 93, 8)),2 => std_logic_vector(to_unsigned( 38, 8)),3 => std_logic_vector(to_unsigned( 29, 8)),4 => std_logic_vector(to_unsigned( 60, 8)),5 => std_logic_vector(to_unsigned( 98, 8)),6 => std_logic_vector(to_unsigned( 24, 8)),7 => std_logic_vector(to_unsigned( 112, 8)),8 => std_logic_vector(to_unsigned( 52, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 61) then
				RAM <= (0 => std_logic_vector(to_unsigned( 94, 8)),1 => std_logic_vector(to_unsigned( 99, 8)),2 => std_logic_vector(to_unsigned( 28, 8)),3 => std_logic_vector(to_unsigned( 77, 8)),4 => std_logic_vector(to_unsigned( 39, 8)),5 => std_logic_vector(to_unsigned( 35, 8)),6 => std_logic_vector(to_unsigned( 83, 8)),7 => std_logic_vector(to_unsigned( 104, 8)),8 => std_logic_vector(to_unsigned( 44, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 62) then
				RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),1 => std_logic_vector(to_unsigned( 111, 8)),2 => std_logic_vector(to_unsigned( 96, 8)),3 => std_logic_vector(to_unsigned( 18, 8)),4 => std_logic_vector(to_unsigned( 23, 8)),5 => std_logic_vector(to_unsigned( 100, 8)),6 => std_logic_vector(to_unsigned( 3, 8)),7 => std_logic_vector(to_unsigned( 30, 8)),8 => std_logic_vector(to_unsigned( 90, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 63) then
				RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),1 => std_logic_vector(to_unsigned( 56, 8)),2 => std_logic_vector(to_unsigned( 32, 8)),3 => std_logic_vector(to_unsigned( 7, 8)),4 => std_logic_vector(to_unsigned( 39, 8)),5 => std_logic_vector(to_unsigned( 52, 8)),6 => std_logic_vector(to_unsigned( 15, 8)),7 => std_logic_vector(to_unsigned( 43, 8)),8 => std_logic_vector(to_unsigned( 0, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 64) then
				RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),1 => std_logic_vector(to_unsigned( 95, 8)),2 => std_logic_vector(to_unsigned( 82, 8)),3 => std_logic_vector(to_unsigned( 51, 8)),4 => std_logic_vector(to_unsigned( 35, 8)),5 => std_logic_vector(to_unsigned( 111, 8)),6 => std_logic_vector(to_unsigned( 117, 8)),7 => std_logic_vector(to_unsigned( 73, 8)),8 => std_logic_vector(to_unsigned( 25, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 65) then
				RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),1 => std_logic_vector(to_unsigned( 43, 8)),2 => std_logic_vector(to_unsigned( 119, 8)),3 => std_logic_vector(to_unsigned( 67, 8)),4 => std_logic_vector(to_unsigned( 47, 8)),5 => std_logic_vector(to_unsigned( 83, 8)),6 => std_logic_vector(to_unsigned( 95, 8)),7 => std_logic_vector(to_unsigned( 22, 8)),8 => std_logic_vector(to_unsigned( 115, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 66) then
				RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),1 => std_logic_vector(to_unsigned( 28, 8)),2 => std_logic_vector(to_unsigned( 95, 8)),3 => std_logic_vector(to_unsigned( 86, 8)),4 => std_logic_vector(to_unsigned( 33, 8)),5 => std_logic_vector(to_unsigned( 110, 8)),6 => std_logic_vector(to_unsigned( 21, 8)),7 => std_logic_vector(to_unsigned( 46, 8)),8 => std_logic_vector(to_unsigned( 62, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 67) then
				RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),1 => std_logic_vector(to_unsigned( 24, 8)),2 => std_logic_vector(to_unsigned( 89, 8)),3 => std_logic_vector(to_unsigned( 94, 8)),4 => std_logic_vector(to_unsigned( 36, 8)),5 => std_logic_vector(to_unsigned( 7, 8)),6 => std_logic_vector(to_unsigned( 50, 8)),7 => std_logic_vector(to_unsigned( 112, 8)),8 => std_logic_vector(to_unsigned( 4, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 68) then
				RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),1 => std_logic_vector(to_unsigned( 15, 8)),2 => std_logic_vector(to_unsigned( 72, 8)),3 => std_logic_vector(to_unsigned( 39, 8)),4 => std_logic_vector(to_unsigned( 104, 8)),5 => std_logic_vector(to_unsigned( 19, 8)),6 => std_logic_vector(to_unsigned( 32, 8)),7 => std_logic_vector(to_unsigned( 9, 8)),8 => std_logic_vector(to_unsigned( 29, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 69) then
				RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),1 => std_logic_vector(to_unsigned( 2, 8)),2 => std_logic_vector(to_unsigned( 17, 8)),3 => std_logic_vector(to_unsigned( 70, 8)),4 => std_logic_vector(to_unsigned( 101, 8)),5 => std_logic_vector(to_unsigned( 46, 8)),6 => std_logic_vector(to_unsigned( 120, 8)),7 => std_logic_vector(to_unsigned( 86, 8)),8 => std_logic_vector(to_unsigned( 82, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 70) then
				RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 77, 8)),3 => std_logic_vector(to_unsigned( 17, 8)),4 => std_logic_vector(to_unsigned( 48, 8)),5 => std_logic_vector(to_unsigned( 56, 8)),6 => std_logic_vector(to_unsigned( 89, 8)),7 => std_logic_vector(to_unsigned( 27, 8)),8 => std_logic_vector(to_unsigned( 125, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 71) then
				RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),1 => std_logic_vector(to_unsigned( 9, 8)),2 => std_logic_vector(to_unsigned( 97, 8)),3 => std_logic_vector(to_unsigned( 63, 8)),4 => std_logic_vector(to_unsigned( 108, 8)),5 => std_logic_vector(to_unsigned( 115, 8)),6 => std_logic_vector(to_unsigned( 83, 8)),7 => std_logic_vector(to_unsigned( 59, 8)),8 => std_logic_vector(to_unsigned( 98, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 72) then
				RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),1 => std_logic_vector(to_unsigned( 76, 8)),2 => std_logic_vector(to_unsigned( 57, 8)),3 => std_logic_vector(to_unsigned( 24, 8)),4 => std_logic_vector(to_unsigned( 115, 8)),5 => std_logic_vector(to_unsigned( 36, 8)),6 => std_logic_vector(to_unsigned( 69, 8)),7 => std_logic_vector(to_unsigned( 64, 8)),8 => std_logic_vector(to_unsigned( 7, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 73) then
				RAM <= (0 => std_logic_vector(to_unsigned( 46, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 21, 8)),3 => std_logic_vector(to_unsigned( 8, 8)),4 => std_logic_vector(to_unsigned( 66, 8)),5 => std_logic_vector(to_unsigned( 58, 8)),6 => std_logic_vector(to_unsigned( 86, 8)),7 => std_logic_vector(to_unsigned( 17, 8)),8 => std_logic_vector(to_unsigned( 37, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 74) then
				RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),1 => std_logic_vector(to_unsigned( 35, 8)),2 => std_logic_vector(to_unsigned( 123, 8)),3 => std_logic_vector(to_unsigned( 40, 8)),4 => std_logic_vector(to_unsigned( 109, 8)),5 => std_logic_vector(to_unsigned( 103, 8)),6 => std_logic_vector(to_unsigned( 44, 8)),7 => std_logic_vector(to_unsigned( 86, 8)),8 => std_logic_vector(to_unsigned( 69, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 75) then
				RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),1 => std_logic_vector(to_unsigned( 86, 8)),2 => std_logic_vector(to_unsigned( 23, 8)),3 => std_logic_vector(to_unsigned( 121, 8)),4 => std_logic_vector(to_unsigned( 109, 8)),5 => std_logic_vector(to_unsigned( 72, 8)),6 => std_logic_vector(to_unsigned( 34, 8)),7 => std_logic_vector(to_unsigned( 113, 8)),8 => std_logic_vector(to_unsigned( 18, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 76) then
				RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),1 => std_logic_vector(to_unsigned( 79, 8)),2 => std_logic_vector(to_unsigned( 72, 8)),3 => std_logic_vector(to_unsigned( 6, 8)),4 => std_logic_vector(to_unsigned( 2, 8)),5 => std_logic_vector(to_unsigned( 102, 8)),6 => std_logic_vector(to_unsigned( 93, 8)),7 => std_logic_vector(to_unsigned( 83, 8)),8 => std_logic_vector(to_unsigned( 88, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 77) then
				RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),1 => std_logic_vector(to_unsigned( 119, 8)),2 => std_logic_vector(to_unsigned( 11, 8)),3 => std_logic_vector(to_unsigned( 68, 8)),4 => std_logic_vector(to_unsigned( 90, 8)),5 => std_logic_vector(to_unsigned( 104, 8)),6 => std_logic_vector(to_unsigned( 109, 8)),7 => std_logic_vector(to_unsigned( 49, 8)),8 => std_logic_vector(to_unsigned( 58, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 78) then
				RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),1 => std_logic_vector(to_unsigned( 27, 8)),2 => std_logic_vector(to_unsigned( 2, 8)),3 => std_logic_vector(to_unsigned( 96, 8)),4 => std_logic_vector(to_unsigned( 108, 8)),5 => std_logic_vector(to_unsigned( 36, 8)),6 => std_logic_vector(to_unsigned( 73, 8)),7 => std_logic_vector(to_unsigned( 7, 8)),8 => std_logic_vector(to_unsigned( 96, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 79) then
				RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),1 => std_logic_vector(to_unsigned( 94, 8)),2 => std_logic_vector(to_unsigned( 85, 8)),3 => std_logic_vector(to_unsigned( 52, 8)),4 => std_logic_vector(to_unsigned( 75, 8)),5 => std_logic_vector(to_unsigned( 29, 8)),6 => std_logic_vector(to_unsigned( 67, 8)),7 => std_logic_vector(to_unsigned( 7, 8)),8 => std_logic_vector(to_unsigned( 112, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 80) then
				RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),1 => std_logic_vector(to_unsigned( 43, 8)),2 => std_logic_vector(to_unsigned( 19, 8)),3 => std_logic_vector(to_unsigned( 66, 8)),4 => std_logic_vector(to_unsigned( 58, 8)),5 => std_logic_vector(to_unsigned( 83, 8)),6 => std_logic_vector(to_unsigned( 118, 8)),7 => std_logic_vector(to_unsigned( 38, 8)),8 => std_logic_vector(to_unsigned( 27, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 81) then
				RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),1 => std_logic_vector(to_unsigned( 12, 8)),2 => std_logic_vector(to_unsigned( 40, 8)),3 => std_logic_vector(to_unsigned( 72, 8)),4 => std_logic_vector(to_unsigned( 111, 8)),5 => std_logic_vector(to_unsigned( 104, 8)),6 => std_logic_vector(to_unsigned( 68, 8)),7 => std_logic_vector(to_unsigned( 16, 8)),8 => std_logic_vector(to_unsigned( 24, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 82) then
				RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),1 => std_logic_vector(to_unsigned( 103, 8)),2 => std_logic_vector(to_unsigned( 95, 8)),3 => std_logic_vector(to_unsigned( 52, 8)),4 => std_logic_vector(to_unsigned( 117, 8)),5 => std_logic_vector(to_unsigned( 81, 8)),6 => std_logic_vector(to_unsigned( 27, 8)),7 => std_logic_vector(to_unsigned( 20, 8)),8 => std_logic_vector(to_unsigned( 90, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 83) then
				RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),1 => std_logic_vector(to_unsigned( 5, 8)),2 => std_logic_vector(to_unsigned( 24, 8)),3 => std_logic_vector(to_unsigned( 31, 8)),4 => std_logic_vector(to_unsigned( 65, 8)),5 => std_logic_vector(to_unsigned( 112, 8)),6 => std_logic_vector(to_unsigned( 90, 8)),7 => std_logic_vector(to_unsigned( 37, 8)),8 => std_logic_vector(to_unsigned( 56, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 84) then
				RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),1 => std_logic_vector(to_unsigned( 63, 8)),2 => std_logic_vector(to_unsigned( 96, 8)),3 => std_logic_vector(to_unsigned( 81, 8)),4 => std_logic_vector(to_unsigned( 116, 8)),5 => std_logic_vector(to_unsigned( 20, 8)),6 => std_logic_vector(to_unsigned( 16, 8)),7 => std_logic_vector(to_unsigned( 12, 8)),8 => std_logic_vector(to_unsigned( 20, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 85) then
				RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),1 => std_logic_vector(to_unsigned( 108, 8)),2 => std_logic_vector(to_unsigned( 78, 8)),3 => std_logic_vector(to_unsigned( 113, 8)),4 => std_logic_vector(to_unsigned( 74, 8)),5 => std_logic_vector(to_unsigned( 7, 8)),6 => std_logic_vector(to_unsigned( 92, 8)),7 => std_logic_vector(to_unsigned( 101, 8)),8 => std_logic_vector(to_unsigned( 93, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 86) then
				RAM <= (0 => std_logic_vector(to_unsigned( 90, 8)),1 => std_logic_vector(to_unsigned( 26, 8)),2 => std_logic_vector(to_unsigned( 124, 8)),3 => std_logic_vector(to_unsigned( 108, 8)),4 => std_logic_vector(to_unsigned( 56, 8)),5 => std_logic_vector(to_unsigned( 36, 8)),6 => std_logic_vector(to_unsigned( 64, 8)),7 => std_logic_vector(to_unsigned( 73, 8)),8 => std_logic_vector(to_unsigned( 31, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 87) then
				RAM <= (0 => std_logic_vector(to_unsigned( 4, 8)),1 => std_logic_vector(to_unsigned( 13, 8)),2 => std_logic_vector(to_unsigned( 67, 8)),3 => std_logic_vector(to_unsigned( 8, 8)),4 => std_logic_vector(to_unsigned( 96, 8)),5 => std_logic_vector(to_unsigned( 88, 8)),6 => std_logic_vector(to_unsigned( 33, 8)),7 => std_logic_vector(to_unsigned( 38, 8)),8 => std_logic_vector(to_unsigned( 121, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 88) then
				RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),1 => std_logic_vector(to_unsigned( 101, 8)),2 => std_logic_vector(to_unsigned( 36, 8)),3 => std_logic_vector(to_unsigned( 4, 8)),4 => std_logic_vector(to_unsigned( 90, 8)),5 => std_logic_vector(to_unsigned( 113, 8)),6 => std_logic_vector(to_unsigned( 45, 8)),7 => std_logic_vector(to_unsigned( 83, 8)),8 => std_logic_vector(to_unsigned( 60, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 89) then
				RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),1 => std_logic_vector(to_unsigned( 63, 8)),2 => std_logic_vector(to_unsigned( 70, 8)),3 => std_logic_vector(to_unsigned( 83, 8)),4 => std_logic_vector(to_unsigned( 99, 8)),5 => std_logic_vector(to_unsigned( 37, 8)),6 => std_logic_vector(to_unsigned( 104, 8)),7 => std_logic_vector(to_unsigned( 55, 8)),8 => std_logic_vector(to_unsigned( 56, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 90) then
				RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),1 => std_logic_vector(to_unsigned( 46, 8)),2 => std_logic_vector(to_unsigned( 96, 8)),3 => std_logic_vector(to_unsigned( 86, 8)),4 => std_logic_vector(to_unsigned( 67, 8)),5 => std_logic_vector(to_unsigned( 63, 8)),6 => std_logic_vector(to_unsigned( 4, 8)),7 => std_logic_vector(to_unsigned( 73, 8)),8 => std_logic_vector(to_unsigned( 112, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 91) then
				RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),1 => std_logic_vector(to_unsigned( 64, 8)),2 => std_logic_vector(to_unsigned( 36, 8)),3 => std_logic_vector(to_unsigned( 120, 8)),4 => std_logic_vector(to_unsigned( 57, 8)),5 => std_logic_vector(to_unsigned( 85, 8)),6 => std_logic_vector(to_unsigned( 94, 8)),7 => std_logic_vector(to_unsigned( 72, 8)),8 => std_logic_vector(to_unsigned( 68, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 92) then
				RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),1 => std_logic_vector(to_unsigned( 65, 8)),2 => std_logic_vector(to_unsigned( 114, 8)),3 => std_logic_vector(to_unsigned( 55, 8)),4 => std_logic_vector(to_unsigned( 92, 8)),5 => std_logic_vector(to_unsigned( 84, 8)),6 => std_logic_vector(to_unsigned( 34, 8)),7 => std_logic_vector(to_unsigned( 11, 8)),8 => std_logic_vector(to_unsigned( 99, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 93) then
				RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),1 => std_logic_vector(to_unsigned( 85, 8)),2 => std_logic_vector(to_unsigned( 116, 8)),3 => std_logic_vector(to_unsigned( 11, 8)),4 => std_logic_vector(to_unsigned( 30, 8)),5 => std_logic_vector(to_unsigned( 43, 8)),6 => std_logic_vector(to_unsigned( 104, 8)),7 => std_logic_vector(to_unsigned( 19, 8)),8 => std_logic_vector(to_unsigned( 37, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 94) then
				RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),1 => std_logic_vector(to_unsigned( 14, 8)),2 => std_logic_vector(to_unsigned( 34, 8)),3 => std_logic_vector(to_unsigned( 72, 8)),4 => std_logic_vector(to_unsigned( 42, 8)),5 => std_logic_vector(to_unsigned( 99, 8)),6 => std_logic_vector(to_unsigned( 6, 8)),7 => std_logic_vector(to_unsigned( 117, 8)),8 => std_logic_vector(to_unsigned( 27, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 95) then
				RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),1 => std_logic_vector(to_unsigned( 122, 8)),2 => std_logic_vector(to_unsigned( 86, 8)),3 => std_logic_vector(to_unsigned( 77, 8)),4 => std_logic_vector(to_unsigned( 19, 8)),5 => std_logic_vector(to_unsigned( 12, 8)),6 => std_logic_vector(to_unsigned( 113, 8)),7 => std_logic_vector(to_unsigned( 52, 8)),8 => std_logic_vector(to_unsigned( 30, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 96) then
				RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),1 => std_logic_vector(to_unsigned( 119, 8)),2 => std_logic_vector(to_unsigned( 107, 8)),3 => std_logic_vector(to_unsigned( 101, 8)),4 => std_logic_vector(to_unsigned( 60, 8)),5 => std_logic_vector(to_unsigned( 113, 8)),6 => std_logic_vector(to_unsigned( 30, 8)),7 => std_logic_vector(to_unsigned( 51, 8)),8 => std_logic_vector(to_unsigned( 50, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 97) then
				RAM <= (0 => std_logic_vector(to_unsigned( 83, 8)),1 => std_logic_vector(to_unsigned( 103, 8)),2 => std_logic_vector(to_unsigned( 75, 8)),3 => std_logic_vector(to_unsigned( 22, 8)),4 => std_logic_vector(to_unsigned( 89, 8)),5 => std_logic_vector(to_unsigned( 96, 8)),6 => std_logic_vector(to_unsigned( 18, 8)),7 => std_logic_vector(to_unsigned( 112, 8)),8 => std_logic_vector(to_unsigned( 82, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 98) then
				RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),1 => std_logic_vector(to_unsigned( 4, 8)),2 => std_logic_vector(to_unsigned( 112, 8)),3 => std_logic_vector(to_unsigned( 33, 8)),4 => std_logic_vector(to_unsigned( 83, 8)),5 => std_logic_vector(to_unsigned( 14, 8)),6 => std_logic_vector(to_unsigned( 44, 8)),7 => std_logic_vector(to_unsigned( 123, 8)),8 => std_logic_vector(to_unsigned( 112, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 99) then
				RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),1 => std_logic_vector(to_unsigned( 39, 8)),2 => std_logic_vector(to_unsigned( 25, 8)),3 => std_logic_vector(to_unsigned( 62, 8)),4 => std_logic_vector(to_unsigned( 3, 8)),5 => std_logic_vector(to_unsigned( 80, 8)),6 => std_logic_vector(to_unsigned( 109, 8)),7 => std_logic_vector(to_unsigned( 44, 8)),8 => std_logic_vector(to_unsigned( 77, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 100) then
				RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),1 => std_logic_vector(to_unsigned( 8, 8)),2 => std_logic_vector(to_unsigned( 28, 8)),3 => std_logic_vector(to_unsigned( 72, 8)),4 => std_logic_vector(to_unsigned( 67, 8)),5 => std_logic_vector(to_unsigned( 87, 8)),6 => std_logic_vector(to_unsigned( 101, 8)),7 => std_logic_vector(to_unsigned( 22, 8)),8 => std_logic_vector(to_unsigned( 2, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 101) then
				RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 5, 8)),3 => std_logic_vector(to_unsigned( 43, 8)),4 => std_logic_vector(to_unsigned( 121, 8)),5 => std_logic_vector(to_unsigned( 78, 8)),6 => std_logic_vector(to_unsigned( 47, 8)),7 => std_logic_vector(to_unsigned( 27, 8)),8 => std_logic_vector(to_unsigned( 19, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 102) then
				RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),1 => std_logic_vector(to_unsigned( 34, 8)),2 => std_logic_vector(to_unsigned( 76, 8)),3 => std_logic_vector(to_unsigned( 3, 8)),4 => std_logic_vector(to_unsigned( 42, 8)),5 => std_logic_vector(to_unsigned( 57, 8)),6 => std_logic_vector(to_unsigned( 18, 8)),7 => std_logic_vector(to_unsigned( 87, 8)),8 => std_logic_vector(to_unsigned( 57, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 103) then
				RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),1 => std_logic_vector(to_unsigned( 86, 8)),2 => std_logic_vector(to_unsigned( 54, 8)),3 => std_logic_vector(to_unsigned( 122, 8)),4 => std_logic_vector(to_unsigned( 2, 8)),5 => std_logic_vector(to_unsigned( 95, 8)),6 => std_logic_vector(to_unsigned( 100, 8)),7 => std_logic_vector(to_unsigned( 48, 8)),8 => std_logic_vector(to_unsigned( 72, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 104) then
				RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),1 => std_logic_vector(to_unsigned( 111, 8)),2 => std_logic_vector(to_unsigned( 38, 8)),3 => std_logic_vector(to_unsigned( 24, 8)),4 => std_logic_vector(to_unsigned( 78, 8)),5 => std_logic_vector(to_unsigned( 58, 8)),6 => std_logic_vector(to_unsigned( 44, 8)),7 => std_logic_vector(to_unsigned( 18, 8)),8 => std_logic_vector(to_unsigned( 17, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 105) then
				RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),1 => std_logic_vector(to_unsigned( 115, 8)),2 => std_logic_vector(to_unsigned( 20, 8)),3 => std_logic_vector(to_unsigned( 44, 8)),4 => std_logic_vector(to_unsigned( 14, 8)),5 => std_logic_vector(to_unsigned( 7, 8)),6 => std_logic_vector(to_unsigned( 121, 8)),7 => std_logic_vector(to_unsigned( 59, 8)),8 => std_logic_vector(to_unsigned( 58, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 106) then
				RAM <= (0 => std_logic_vector(to_unsigned( 53, 8)),1 => std_logic_vector(to_unsigned( 84, 8)),2 => std_logic_vector(to_unsigned( 4, 8)),3 => std_logic_vector(to_unsigned( 94, 8)),4 => std_logic_vector(to_unsigned( 17, 8)),5 => std_logic_vector(to_unsigned( 22, 8)),6 => std_logic_vector(to_unsigned( 98, 8)),7 => std_logic_vector(to_unsigned( 42, 8)),8 => std_logic_vector(to_unsigned( 109, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 107) then
				RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),1 => std_logic_vector(to_unsigned( 53, 8)),2 => std_logic_vector(to_unsigned( 66, 8)),3 => std_logic_vector(to_unsigned( 112, 8)),4 => std_logic_vector(to_unsigned( 25, 8)),5 => std_logic_vector(to_unsigned( 3, 8)),6 => std_logic_vector(to_unsigned( 89, 8)),7 => std_logic_vector(to_unsigned( 117, 8)),8 => std_logic_vector(to_unsigned( 69, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 108) then
				RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),1 => std_logic_vector(to_unsigned( 1, 8)),2 => std_logic_vector(to_unsigned( 46, 8)),3 => std_logic_vector(to_unsigned( 35, 8)),4 => std_logic_vector(to_unsigned( 29, 8)),5 => std_logic_vector(to_unsigned( 41, 8)),6 => std_logic_vector(to_unsigned( 104, 8)),7 => std_logic_vector(to_unsigned( 23, 8)),8 => std_logic_vector(to_unsigned( 7, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 109) then
				RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),1 => std_logic_vector(to_unsigned( 14, 8)),2 => std_logic_vector(to_unsigned( 80, 8)),3 => std_logic_vector(to_unsigned( 1, 8)),4 => std_logic_vector(to_unsigned( 44, 8)),5 => std_logic_vector(to_unsigned( 30, 8)),6 => std_logic_vector(to_unsigned( 70, 8)),7 => std_logic_vector(to_unsigned( 96, 8)),8 => std_logic_vector(to_unsigned( 89, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 110) then
				RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),1 => std_logic_vector(to_unsigned( 124, 8)),2 => std_logic_vector(to_unsigned( 15, 8)),3 => std_logic_vector(to_unsigned( 75, 8)),4 => std_logic_vector(to_unsigned( 63, 8)),5 => std_logic_vector(to_unsigned( 106, 8)),6 => std_logic_vector(to_unsigned( 56, 8)),7 => std_logic_vector(to_unsigned( 81, 8)),8 => std_logic_vector(to_unsigned( 16, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 111) then
				RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),1 => std_logic_vector(to_unsigned( 102, 8)),2 => std_logic_vector(to_unsigned( 9, 8)),3 => std_logic_vector(to_unsigned( 121, 8)),4 => std_logic_vector(to_unsigned( 27, 8)),5 => std_logic_vector(to_unsigned( 20, 8)),6 => std_logic_vector(to_unsigned( 111, 8)),7 => std_logic_vector(to_unsigned( 80, 8)),8 => std_logic_vector(to_unsigned( 88, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 112) then
				RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),1 => std_logic_vector(to_unsigned( 99, 8)),2 => std_logic_vector(to_unsigned( 44, 8)),3 => std_logic_vector(to_unsigned( 50, 8)),4 => std_logic_vector(to_unsigned( 121, 8)),5 => std_logic_vector(to_unsigned( 70, 8)),6 => std_logic_vector(to_unsigned( 113, 8)),7 => std_logic_vector(to_unsigned( 34, 8)),8 => std_logic_vector(to_unsigned( 114, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 113) then
				RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),1 => std_logic_vector(to_unsigned( 94, 8)),2 => std_logic_vector(to_unsigned( 52, 8)),3 => std_logic_vector(to_unsigned( 27, 8)),4 => std_logic_vector(to_unsigned( 39, 8)),5 => std_logic_vector(to_unsigned( 60, 8)),6 => std_logic_vector(to_unsigned( 114, 8)),7 => std_logic_vector(to_unsigned( 77, 8)),8 => std_logic_vector(to_unsigned( 11, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 114) then
				RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),1 => std_logic_vector(to_unsigned( 48, 8)),2 => std_logic_vector(to_unsigned( 96, 8)),3 => std_logic_vector(to_unsigned( 102, 8)),4 => std_logic_vector(to_unsigned( 64, 8)),5 => std_logic_vector(to_unsigned( 113, 8)),6 => std_logic_vector(to_unsigned( 109, 8)),7 => std_logic_vector(to_unsigned( 56, 8)),8 => std_logic_vector(to_unsigned( 55, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 115) then
				RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),1 => std_logic_vector(to_unsigned( 89, 8)),2 => std_logic_vector(to_unsigned( 94, 8)),3 => std_logic_vector(to_unsigned( 120, 8)),4 => std_logic_vector(to_unsigned( 57, 8)),5 => std_logic_vector(to_unsigned( 110, 8)),6 => std_logic_vector(to_unsigned( 31, 8)),7 => std_logic_vector(to_unsigned( 63, 8)),8 => std_logic_vector(to_unsigned( 10, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 116) then
				RAM <= (0 => std_logic_vector(to_unsigned( 8, 8)),1 => std_logic_vector(to_unsigned( 99, 8)),2 => std_logic_vector(to_unsigned( 30, 8)),3 => std_logic_vector(to_unsigned( 85, 8)),4 => std_logic_vector(to_unsigned( 109, 8)),5 => std_logic_vector(to_unsigned( 55, 8)),6 => std_logic_vector(to_unsigned( 23, 8)),7 => std_logic_vector(to_unsigned( 16, 8)),8 => std_logic_vector(to_unsigned( 3, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 117) then
				RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),1 => std_logic_vector(to_unsigned( 49, 8)),2 => std_logic_vector(to_unsigned( 110, 8)),3 => std_logic_vector(to_unsigned( 81, 8)),4 => std_logic_vector(to_unsigned( 121, 8)),5 => std_logic_vector(to_unsigned( 31, 8)),6 => std_logic_vector(to_unsigned( 53, 8)),7 => std_logic_vector(to_unsigned( 25, 8)),8 => std_logic_vector(to_unsigned( 57, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 118) then
				RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),1 => std_logic_vector(to_unsigned( 17, 8)),2 => std_logic_vector(to_unsigned( 90, 8)),3 => std_logic_vector(to_unsigned( 79, 8)),4 => std_logic_vector(to_unsigned( 41, 8)),5 => std_logic_vector(to_unsigned( 116, 8)),6 => std_logic_vector(to_unsigned( 55, 8)),7 => std_logic_vector(to_unsigned( 66, 8)),8 => std_logic_vector(to_unsigned( 64, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 119) then
				RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),1 => std_logic_vector(to_unsigned( 14, 8)),2 => std_logic_vector(to_unsigned( 82, 8)),3 => std_logic_vector(to_unsigned( 7, 8)),4 => std_logic_vector(to_unsigned( 72, 8)),5 => std_logic_vector(to_unsigned( 36, 8)),6 => std_logic_vector(to_unsigned( 41, 8)),7 => std_logic_vector(to_unsigned( 57, 8)),8 => std_logic_vector(to_unsigned( 13, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 120) then
				RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),1 => std_logic_vector(to_unsigned( 83, 8)),2 => std_logic_vector(to_unsigned( 16, 8)),3 => std_logic_vector(to_unsigned( 114, 8)),4 => std_logic_vector(to_unsigned( 45, 8)),5 => std_logic_vector(to_unsigned( 22, 8)),6 => std_logic_vector(to_unsigned( 93, 8)),7 => std_logic_vector(to_unsigned( 55, 8)),8 => std_logic_vector(to_unsigned( 27, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 121) then
				RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),1 => std_logic_vector(to_unsigned( 121, 8)),2 => std_logic_vector(to_unsigned( 86, 8)),3 => std_logic_vector(to_unsigned( 98, 8)),4 => std_logic_vector(to_unsigned( 7, 8)),5 => std_logic_vector(to_unsigned( 24, 8)),6 => std_logic_vector(to_unsigned( 2, 8)),7 => std_logic_vector(to_unsigned( 70, 8)),8 => std_logic_vector(to_unsigned( 74, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 122) then
				RAM <= (0 => std_logic_vector(to_unsigned( 77, 8)),1 => std_logic_vector(to_unsigned( 14, 8)),2 => std_logic_vector(to_unsigned( 28, 8)),3 => std_logic_vector(to_unsigned( 106, 8)),4 => std_logic_vector(to_unsigned( 19, 8)),5 => std_logic_vector(to_unsigned( 85, 8)),6 => std_logic_vector(to_unsigned( 36, 8)),7 => std_logic_vector(to_unsigned( 51, 8)),8 => std_logic_vector(to_unsigned( 19, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 123) then
				RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),1 => std_logic_vector(to_unsigned( 77, 8)),2 => std_logic_vector(to_unsigned( 111, 8)),3 => std_logic_vector(to_unsigned( 93, 8)),4 => std_logic_vector(to_unsigned( 85, 8)),5 => std_logic_vector(to_unsigned( 4, 8)),6 => std_logic_vector(to_unsigned( 68, 8)),7 => std_logic_vector(to_unsigned( 33, 8)),8 => std_logic_vector(to_unsigned( 72, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 124) then
				RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),1 => std_logic_vector(to_unsigned( 111, 8)),2 => std_logic_vector(to_unsigned( 16, 8)),3 => std_logic_vector(to_unsigned( 29, 8)),4 => std_logic_vector(to_unsigned( 22, 8)),5 => std_logic_vector(to_unsigned( 35, 8)),6 => std_logic_vector(to_unsigned( 55, 8)),7 => std_logic_vector(to_unsigned( 70, 8)),8 => std_logic_vector(to_unsigned( 83, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 125) then
				RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),1 => std_logic_vector(to_unsigned( 4, 8)),2 => std_logic_vector(to_unsigned( 97, 8)),3 => std_logic_vector(to_unsigned( 43, 8)),4 => std_logic_vector(to_unsigned( 88, 8)),5 => std_logic_vector(to_unsigned( 21, 8)),6 => std_logic_vector(to_unsigned( 54, 8)),7 => std_logic_vector(to_unsigned( 107, 8)),8 => std_logic_vector(to_unsigned( 55, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 126) then
				RAM <= (0 => std_logic_vector(to_unsigned( 90, 8)),1 => std_logic_vector(to_unsigned( 27, 8)),2 => std_logic_vector(to_unsigned( 35, 8)),3 => std_logic_vector(to_unsigned( 82, 8)),4 => std_logic_vector(to_unsigned( 98, 8)),5 => std_logic_vector(to_unsigned( 16, 8)),6 => std_logic_vector(to_unsigned( 68, 8)),7 => std_logic_vector(to_unsigned( 7, 8)),8 => std_logic_vector(to_unsigned( 48, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 127) then
				RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),1 => std_logic_vector(to_unsigned( 81, 8)),2 => std_logic_vector(to_unsigned( 102, 8)),3 => std_logic_vector(to_unsigned( 70, 8)),4 => std_logic_vector(to_unsigned( 96, 8)),5 => std_logic_vector(to_unsigned( 29, 8)),6 => std_logic_vector(to_unsigned( 58, 8)),7 => std_logic_vector(to_unsigned( 92, 8)),8 => std_logic_vector(to_unsigned( 41, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 128) then
				RAM <= (0 => std_logic_vector(to_unsigned( 70, 8)),1 => std_logic_vector(to_unsigned( 77, 8)),2 => std_logic_vector(to_unsigned( 40, 8)),3 => std_logic_vector(to_unsigned( 111, 8)),4 => std_logic_vector(to_unsigned( 36, 8)),5 => std_logic_vector(to_unsigned( 87, 8)),6 => std_logic_vector(to_unsigned( 6, 8)),7 => std_logic_vector(to_unsigned( 29, 8)),8 => std_logic_vector(to_unsigned( 17, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 129) then
				RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),1 => std_logic_vector(to_unsigned( 93, 8)),2 => std_logic_vector(to_unsigned( 124, 8)),3 => std_logic_vector(to_unsigned( 75, 8)),4 => std_logic_vector(to_unsigned( 105, 8)),5 => std_logic_vector(to_unsigned( 2, 8)),6 => std_logic_vector(to_unsigned( 85, 8)),7 => std_logic_vector(to_unsigned( 39, 8)),8 => std_logic_vector(to_unsigned( 5, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 130) then
				RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),1 => std_logic_vector(to_unsigned( 13, 8)),2 => std_logic_vector(to_unsigned( 78, 8)),3 => std_logic_vector(to_unsigned( 61, 8)),4 => std_logic_vector(to_unsigned( 109, 8)),5 => std_logic_vector(to_unsigned( 96, 8)),6 => std_logic_vector(to_unsigned( 85, 8)),7 => std_logic_vector(to_unsigned( 50, 8)),8 => std_logic_vector(to_unsigned( 33, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 131) then
				RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),1 => std_logic_vector(to_unsigned( 14, 8)),2 => std_logic_vector(to_unsigned( 123, 8)),3 => std_logic_vector(to_unsigned( 108, 8)),4 => std_logic_vector(to_unsigned( 1, 8)),5 => std_logic_vector(to_unsigned( 115, 8)),6 => std_logic_vector(to_unsigned( 40, 8)),7 => std_logic_vector(to_unsigned( 9, 8)),8 => std_logic_vector(to_unsigned( 93, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 132) then
				RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),1 => std_logic_vector(to_unsigned( 51, 8)),2 => std_logic_vector(to_unsigned( 55, 8)),3 => std_logic_vector(to_unsigned( 116, 8)),4 => std_logic_vector(to_unsigned( 18, 8)),5 => std_logic_vector(to_unsigned( 66, 8)),6 => std_logic_vector(to_unsigned( 61, 8)),7 => std_logic_vector(to_unsigned( 86, 8)),8 => std_logic_vector(to_unsigned( 17, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 133) then
				RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),1 => std_logic_vector(to_unsigned( 71, 8)),2 => std_logic_vector(to_unsigned( 4, 8)),3 => std_logic_vector(to_unsigned( 16, 8)),4 => std_logic_vector(to_unsigned( 92, 8)),5 => std_logic_vector(to_unsigned( 85, 8)),6 => std_logic_vector(to_unsigned( 51, 8)),7 => std_logic_vector(to_unsigned( 104, 8)),8 => std_logic_vector(to_unsigned( 41, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 134) then
				RAM <= (0 => std_logic_vector(to_unsigned( 84, 8)),1 => std_logic_vector(to_unsigned( 122, 8)),2 => std_logic_vector(to_unsigned( 19, 8)),3 => std_logic_vector(to_unsigned( 52, 8)),4 => std_logic_vector(to_unsigned( 12, 8)),5 => std_logic_vector(to_unsigned( 100, 8)),6 => std_logic_vector(to_unsigned( 32, 8)),7 => std_logic_vector(to_unsigned( 73, 8)),8 => std_logic_vector(to_unsigned( 19, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 135) then
				RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),1 => std_logic_vector(to_unsigned( 65, 8)),2 => std_logic_vector(to_unsigned( 103, 8)),3 => std_logic_vector(to_unsigned( 93, 8)),4 => std_logic_vector(to_unsigned( 34, 8)),5 => std_logic_vector(to_unsigned( 116, 8)),6 => std_logic_vector(to_unsigned( 77, 8)),7 => std_logic_vector(to_unsigned( 124, 8)),8 => std_logic_vector(to_unsigned( 40, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 136) then
				RAM <= (0 => std_logic_vector(to_unsigned( 88, 8)),1 => std_logic_vector(to_unsigned( 80, 8)),2 => std_logic_vector(to_unsigned( 62, 8)),3 => std_logic_vector(to_unsigned( 37, 8)),4 => std_logic_vector(to_unsigned( 54, 8)),5 => std_logic_vector(to_unsigned( 93, 8)),6 => std_logic_vector(to_unsigned( 24, 8)),7 => std_logic_vector(to_unsigned( 1, 8)),8 => std_logic_vector(to_unsigned( 23, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 137) then
				RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),1 => std_logic_vector(to_unsigned( 95, 8)),2 => std_logic_vector(to_unsigned( 27, 8)),3 => std_logic_vector(to_unsigned( 37, 8)),4 => std_logic_vector(to_unsigned( 119, 8)),5 => std_logic_vector(to_unsigned( 64, 8)),6 => std_logic_vector(to_unsigned( 68, 8)),7 => std_logic_vector(to_unsigned( 91, 8)),8 => std_logic_vector(to_unsigned( 31, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 138) then
				RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 19, 8)),3 => std_logic_vector(to_unsigned( 51, 8)),4 => std_logic_vector(to_unsigned( 36, 8)),5 => std_logic_vector(to_unsigned( 29, 8)),6 => std_logic_vector(to_unsigned( 9, 8)),7 => std_logic_vector(to_unsigned( 3, 8)),8 => std_logic_vector(to_unsigned( 96, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 139) then
				RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),1 => std_logic_vector(to_unsigned( 65, 8)),2 => std_logic_vector(to_unsigned( 109, 8)),3 => std_logic_vector(to_unsigned( 99, 8)),4 => std_logic_vector(to_unsigned( 37, 8)),5 => std_logic_vector(to_unsigned( 104, 8)),6 => std_logic_vector(to_unsigned( 51, 8)),7 => std_logic_vector(to_unsigned( 6, 8)),8 => std_logic_vector(to_unsigned( 3, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 140) then
				RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),1 => std_logic_vector(to_unsigned( 20, 8)),2 => std_logic_vector(to_unsigned( 12, 8)),3 => std_logic_vector(to_unsigned( 70, 8)),4 => std_logic_vector(to_unsigned( 59, 8)),5 => std_logic_vector(to_unsigned( 42, 8)),6 => std_logic_vector(to_unsigned( 120, 8)),7 => std_logic_vector(to_unsigned( 111, 8)),8 => std_logic_vector(to_unsigned( 42, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 141) then
				RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),1 => std_logic_vector(to_unsigned( 23, 8)),2 => std_logic_vector(to_unsigned( 28, 8)),3 => std_logic_vector(to_unsigned( 77, 8)),4 => std_logic_vector(to_unsigned( 38, 8)),5 => std_logic_vector(to_unsigned( 52, 8)),6 => std_logic_vector(to_unsigned( 56, 8)),7 => std_logic_vector(to_unsigned( 9, 8)),8 => std_logic_vector(to_unsigned( 112, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 142) then
				RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),1 => std_logic_vector(to_unsigned( 51, 8)),2 => std_logic_vector(to_unsigned( 96, 8)),3 => std_logic_vector(to_unsigned( 0, 8)),4 => std_logic_vector(to_unsigned( 10, 8)),5 => std_logic_vector(to_unsigned( 28, 8)),6 => std_logic_vector(to_unsigned( 47, 8)),7 => std_logic_vector(to_unsigned( 39, 8)),8 => std_logic_vector(to_unsigned( 18, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 143) then
				RAM <= (0 => std_logic_vector(to_unsigned( 62, 8)),1 => std_logic_vector(to_unsigned( 119, 8)),2 => std_logic_vector(to_unsigned( 58, 8)),3 => std_logic_vector(to_unsigned( 32, 8)),4 => std_logic_vector(to_unsigned( 72, 8)),5 => std_logic_vector(to_unsigned( 96, 8)),6 => std_logic_vector(to_unsigned( 0, 8)),7 => std_logic_vector(to_unsigned( 67, 8)),8 => std_logic_vector(to_unsigned( 64, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 144) then
				RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),1 => std_logic_vector(to_unsigned( 41, 8)),2 => std_logic_vector(to_unsigned( 98, 8)),3 => std_logic_vector(to_unsigned( 113, 8)),4 => std_logic_vector(to_unsigned( 58, 8)),5 => std_logic_vector(to_unsigned( 30, 8)),6 => std_logic_vector(to_unsigned( 85, 8)),7 => std_logic_vector(to_unsigned( 37, 8)),8 => std_logic_vector(to_unsigned( 25, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 145) then
				RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),1 => std_logic_vector(to_unsigned( 71, 8)),2 => std_logic_vector(to_unsigned( 109, 8)),3 => std_logic_vector(to_unsigned( 115, 8)),4 => std_logic_vector(to_unsigned( 2, 8)),5 => std_logic_vector(to_unsigned( 59, 8)),6 => std_logic_vector(to_unsigned( 15, 8)),7 => std_logic_vector(to_unsigned( 80, 8)),8 => std_logic_vector(to_unsigned( 40, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 146) then
				RAM <= (0 => std_logic_vector(to_unsigned( 114, 8)),1 => std_logic_vector(to_unsigned( 67, 8)),2 => std_logic_vector(to_unsigned( 22, 8)),3 => std_logic_vector(to_unsigned( 105, 8)),4 => std_logic_vector(to_unsigned( 32, 8)),5 => std_logic_vector(to_unsigned( 57, 8)),6 => std_logic_vector(to_unsigned( 78, 8)),7 => std_logic_vector(to_unsigned( 74, 8)),8 => std_logic_vector(to_unsigned( 56, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 147) then
				RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),1 => std_logic_vector(to_unsigned( 12, 8)),2 => std_logic_vector(to_unsigned( 83, 8)),3 => std_logic_vector(to_unsigned( 24, 8)),4 => std_logic_vector(to_unsigned( 94, 8)),5 => std_logic_vector(to_unsigned( 106, 8)),6 => std_logic_vector(to_unsigned( 115, 8)),7 => std_logic_vector(to_unsigned( 89, 8)),8 => std_logic_vector(to_unsigned( 56, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 148) then
				RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),1 => std_logic_vector(to_unsigned( 98, 8)),2 => std_logic_vector(to_unsigned( 83, 8)),3 => std_logic_vector(to_unsigned( 67, 8)),4 => std_logic_vector(to_unsigned( 122, 8)),5 => std_logic_vector(to_unsigned( 29, 8)),6 => std_logic_vector(to_unsigned( 52, 8)),7 => std_logic_vector(to_unsigned( 37, 8)),8 => std_logic_vector(to_unsigned( 58, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 149) then
				RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),1 => std_logic_vector(to_unsigned( 20, 8)),2 => std_logic_vector(to_unsigned( 80, 8)),3 => std_logic_vector(to_unsigned( 61, 8)),4 => std_logic_vector(to_unsigned( 117, 8)),5 => std_logic_vector(to_unsigned( 89, 8)),6 => std_logic_vector(to_unsigned( 32, 8)),7 => std_logic_vector(to_unsigned( 93, 8)),8 => std_logic_vector(to_unsigned( 89, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 150) then
				RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),1 => std_logic_vector(to_unsigned( 121, 8)),2 => std_logic_vector(to_unsigned( 90, 8)),3 => std_logic_vector(to_unsigned( 49, 8)),4 => std_logic_vector(to_unsigned( 25, 8)),5 => std_logic_vector(to_unsigned( 69, 8)),6 => std_logic_vector(to_unsigned( 0, 8)),7 => std_logic_vector(to_unsigned( 15, 8)),8 => std_logic_vector(to_unsigned( 47, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 151) then
				RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),1 => std_logic_vector(to_unsigned( 111, 8)),2 => std_logic_vector(to_unsigned( 85, 8)),3 => std_logic_vector(to_unsigned( 79, 8)),4 => std_logic_vector(to_unsigned( 2, 8)),5 => std_logic_vector(to_unsigned( 34, 8)),6 => std_logic_vector(to_unsigned( 47, 8)),7 => std_logic_vector(to_unsigned( 105, 8)),8 => std_logic_vector(to_unsigned( 11, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 152) then
				RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),1 => std_logic_vector(to_unsigned( 85, 8)),2 => std_logic_vector(to_unsigned( 3, 8)),3 => std_logic_vector(to_unsigned( 121, 8)),4 => std_logic_vector(to_unsigned( 43, 8)),5 => std_logic_vector(to_unsigned( 76, 8)),6 => std_logic_vector(to_unsigned( 94, 8)),7 => std_logic_vector(to_unsigned( 109, 8)),8 => std_logic_vector(to_unsigned( 21, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 153) then
				RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),1 => std_logic_vector(to_unsigned( 46, 8)),2 => std_logic_vector(to_unsigned( 113, 8)),3 => std_logic_vector(to_unsigned( 106, 8)),4 => std_logic_vector(to_unsigned( 42, 8)),5 => std_logic_vector(to_unsigned( 6, 8)),6 => std_logic_vector(to_unsigned( 89, 8)),7 => std_logic_vector(to_unsigned( 124, 8)),8 => std_logic_vector(to_unsigned( 10, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 154) then
				RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),1 => std_logic_vector(to_unsigned( 109, 8)),2 => std_logic_vector(to_unsigned( 58, 8)),3 => std_logic_vector(to_unsigned( 34, 8)),4 => std_logic_vector(to_unsigned( 64, 8)),5 => std_logic_vector(to_unsigned( 13, 8)),6 => std_logic_vector(to_unsigned( 116, 8)),7 => std_logic_vector(to_unsigned( 73, 8)),8 => std_logic_vector(to_unsigned( 56, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 155) then
				RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),1 => std_logic_vector(to_unsigned( 80, 8)),2 => std_logic_vector(to_unsigned( 57, 8)),3 => std_logic_vector(to_unsigned( 112, 8)),4 => std_logic_vector(to_unsigned( 52, 8)),5 => std_logic_vector(to_unsigned( 96, 8)),6 => std_logic_vector(to_unsigned( 62, 8)),7 => std_logic_vector(to_unsigned( 40, 8)),8 => std_logic_vector(to_unsigned( 49, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 156) then
				RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),1 => std_logic_vector(to_unsigned( 37, 8)),2 => std_logic_vector(to_unsigned( 94, 8)),3 => std_logic_vector(to_unsigned( 27, 8)),4 => std_logic_vector(to_unsigned( 87, 8)),5 => std_logic_vector(to_unsigned( 18, 8)),6 => std_logic_vector(to_unsigned( 64, 8)),7 => std_logic_vector(to_unsigned( 5, 8)),8 => std_logic_vector(to_unsigned( 17, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 157) then
				RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),1 => std_logic_vector(to_unsigned( 9, 8)),2 => std_logic_vector(to_unsigned( 56, 8)),3 => std_logic_vector(to_unsigned( 85, 8)),4 => std_logic_vector(to_unsigned( 99, 8)),5 => std_logic_vector(to_unsigned( 32, 8)),6 => std_logic_vector(to_unsigned( 65, 8)),7 => std_logic_vector(to_unsigned( 1, 8)),8 => std_logic_vector(to_unsigned( 41, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 158) then
				RAM <= (0 => std_logic_vector(to_unsigned( 38, 8)),1 => std_logic_vector(to_unsigned( 5, 8)),2 => std_logic_vector(to_unsigned( 53, 8)),3 => std_logic_vector(to_unsigned( 80, 8)),4 => std_logic_vector(to_unsigned( 44, 8)),5 => std_logic_vector(to_unsigned( 119, 8)),6 => std_logic_vector(to_unsigned( 109, 8)),7 => std_logic_vector(to_unsigned( 10, 8)),8 => std_logic_vector(to_unsigned( 2, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 159) then
				RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),1 => std_logic_vector(to_unsigned( 44, 8)),2 => std_logic_vector(to_unsigned( 23, 8)),3 => std_logic_vector(to_unsigned( 31, 8)),4 => std_logic_vector(to_unsigned( 0, 8)),5 => std_logic_vector(to_unsigned( 62, 8)),6 => std_logic_vector(to_unsigned( 52, 8)),7 => std_logic_vector(to_unsigned( 97, 8)),8 => std_logic_vector(to_unsigned( 61, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 160) then
				RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),1 => std_logic_vector(to_unsigned( 46, 8)),2 => std_logic_vector(to_unsigned( 120, 8)),3 => std_logic_vector(to_unsigned( 5, 8)),4 => std_logic_vector(to_unsigned( 100, 8)),5 => std_logic_vector(to_unsigned( 61, 8)),6 => std_logic_vector(to_unsigned( 107, 8)),7 => std_logic_vector(to_unsigned( 18, 8)),8 => std_logic_vector(to_unsigned( 71, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 161) then
				RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),1 => std_logic_vector(to_unsigned( 22, 8)),2 => std_logic_vector(to_unsigned( 80, 8)),3 => std_logic_vector(to_unsigned( 57, 8)),4 => std_logic_vector(to_unsigned( 14, 8)),5 => std_logic_vector(to_unsigned( 63, 8)),6 => std_logic_vector(to_unsigned( 91, 8)),7 => std_logic_vector(to_unsigned( 114, 8)),8 => std_logic_vector(to_unsigned( 126, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 162) then
				RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),1 => std_logic_vector(to_unsigned( 118, 8)),2 => std_logic_vector(to_unsigned( 5, 8)),3 => std_logic_vector(to_unsigned( 19, 8)),4 => std_logic_vector(to_unsigned( 95, 8)),5 => std_logic_vector(to_unsigned( 10, 8)),6 => std_logic_vector(to_unsigned( 35, 8)),7 => std_logic_vector(to_unsigned( 68, 8)),8 => std_logic_vector(to_unsigned( 33, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 163) then
				RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),1 => std_logic_vector(to_unsigned( 56, 8)),2 => std_logic_vector(to_unsigned( 30, 8)),3 => std_logic_vector(to_unsigned( 3, 8)),4 => std_logic_vector(to_unsigned( 35, 8)),5 => std_logic_vector(to_unsigned( 47, 8)),6 => std_logic_vector(to_unsigned( 119, 8)),7 => std_logic_vector(to_unsigned( 8, 8)),8 => std_logic_vector(to_unsigned( 39, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 164) then
				RAM <= (0 => std_logic_vector(to_unsigned( 39, 8)),1 => std_logic_vector(to_unsigned( 3, 8)),2 => std_logic_vector(to_unsigned( 110, 8)),3 => std_logic_vector(to_unsigned( 14, 8)),4 => std_logic_vector(to_unsigned( 45, 8)),5 => std_logic_vector(to_unsigned( 92, 8)),6 => std_logic_vector(to_unsigned( 26, 8)),7 => std_logic_vector(to_unsigned( 119, 8)),8 => std_logic_vector(to_unsigned( 46, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 165) then
				RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),1 => std_logic_vector(to_unsigned( 84, 8)),2 => std_logic_vector(to_unsigned( 89, 8)),3 => std_logic_vector(to_unsigned( 30, 8)),4 => std_logic_vector(to_unsigned( 76, 8)),5 => std_logic_vector(to_unsigned( 68, 8)),6 => std_logic_vector(to_unsigned( 50, 8)),7 => std_logic_vector(to_unsigned( 36, 8)),8 => std_logic_vector(to_unsigned( 101, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 166) then
				RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),1 => std_logic_vector(to_unsigned( 24, 8)),2 => std_logic_vector(to_unsigned( 121, 8)),3 => std_logic_vector(to_unsigned( 16, 8)),4 => std_logic_vector(to_unsigned( 105, 8)),5 => std_logic_vector(to_unsigned( 50, 8)),6 => std_logic_vector(to_unsigned( 88, 8)),7 => std_logic_vector(to_unsigned( 64, 8)),8 => std_logic_vector(to_unsigned( 95, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 167) then
				RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),1 => std_logic_vector(to_unsigned( 68, 8)),2 => std_logic_vector(to_unsigned( 85, 8)),3 => std_logic_vector(to_unsigned( 26, 8)),4 => std_logic_vector(to_unsigned( 124, 8)),5 => std_logic_vector(to_unsigned( 37, 8)),6 => std_logic_vector(to_unsigned( 22, 8)),7 => std_logic_vector(to_unsigned( 91, 8)),8 => std_logic_vector(to_unsigned( 126, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 168) then
				RAM <= (0 => std_logic_vector(to_unsigned( 114, 8)),1 => std_logic_vector(to_unsigned( 79, 8)),2 => std_logic_vector(to_unsigned( 7, 8)),3 => std_logic_vector(to_unsigned( 106, 8)),4 => std_logic_vector(to_unsigned( 100, 8)),5 => std_logic_vector(to_unsigned( 67, 8)),6 => std_logic_vector(to_unsigned( 91, 8)),7 => std_logic_vector(to_unsigned( 14, 8)),8 => std_logic_vector(to_unsigned( 36, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 169) then
				RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),1 => std_logic_vector(to_unsigned( 17, 8)),2 => std_logic_vector(to_unsigned( 121, 8)),3 => std_logic_vector(to_unsigned( 49, 8)),4 => std_logic_vector(to_unsigned( 90, 8)),5 => std_logic_vector(to_unsigned( 97, 8)),6 => std_logic_vector(to_unsigned( 7, 8)),7 => std_logic_vector(to_unsigned( 78, 8)),8 => std_logic_vector(to_unsigned( 44, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 170) then
				RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),1 => std_logic_vector(to_unsigned( 33, 8)),2 => std_logic_vector(to_unsigned( 124, 8)),3 => std_logic_vector(to_unsigned( 61, 8)),4 => std_logic_vector(to_unsigned( 7, 8)),5 => std_logic_vector(to_unsigned( 95, 8)),6 => std_logic_vector(to_unsigned( 42, 8)),7 => std_logic_vector(to_unsigned( 120, 8)),8 => std_logic_vector(to_unsigned( 77, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 171) then
				RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),1 => std_logic_vector(to_unsigned( 113, 8)),2 => std_logic_vector(to_unsigned( 60, 8)),3 => std_logic_vector(to_unsigned( 87, 8)),4 => std_logic_vector(to_unsigned( 18, 8)),5 => std_logic_vector(to_unsigned( 11, 8)),6 => std_logic_vector(to_unsigned( 103, 8)),7 => std_logic_vector(to_unsigned( 93, 8)),8 => std_logic_vector(to_unsigned( 64, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 172) then
				RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),1 => std_logic_vector(to_unsigned( 10, 8)),2 => std_logic_vector(to_unsigned( 2, 8)),3 => std_logic_vector(to_unsigned( 46, 8)),4 => std_logic_vector(to_unsigned( 111, 8)),5 => std_logic_vector(to_unsigned( 69, 8)),6 => std_logic_vector(to_unsigned( 55, 8)),7 => std_logic_vector(to_unsigned( 19, 8)),8 => std_logic_vector(to_unsigned( 11, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 173) then
				RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),1 => std_logic_vector(to_unsigned( 21, 8)),2 => std_logic_vector(to_unsigned( 2, 8)),3 => std_logic_vector(to_unsigned( 68, 8)),4 => std_logic_vector(to_unsigned( 124, 8)),5 => std_logic_vector(to_unsigned( 37, 8)),6 => std_logic_vector(to_unsigned( 84, 8)),7 => std_logic_vector(to_unsigned( 64, 8)),8 => std_logic_vector(to_unsigned( 90, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 174) then
				RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),1 => std_logic_vector(to_unsigned( 29, 8)),2 => std_logic_vector(to_unsigned( 1, 8)),3 => std_logic_vector(to_unsigned( 113, 8)),4 => std_logic_vector(to_unsigned( 93, 8)),5 => std_logic_vector(to_unsigned( 84, 8)),6 => std_logic_vector(to_unsigned( 34, 8)),7 => std_logic_vector(to_unsigned( 102, 8)),8 => std_logic_vector(to_unsigned( 35, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 175) then
				RAM <= (0 => std_logic_vector(to_unsigned( 115, 8)),1 => std_logic_vector(to_unsigned( 40, 8)),2 => std_logic_vector(to_unsigned( 71, 8)),3 => std_logic_vector(to_unsigned( 33, 8)),4 => std_logic_vector(to_unsigned( 45, 8)),5 => std_logic_vector(to_unsigned( 8, 8)),6 => std_logic_vector(to_unsigned( 27, 8)),7 => std_logic_vector(to_unsigned( 20, 8)),8 => std_logic_vector(to_unsigned( 97, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 176) then
				RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),1 => std_logic_vector(to_unsigned( 74, 8)),2 => std_logic_vector(to_unsigned( 99, 8)),3 => std_logic_vector(to_unsigned( 59, 8)),4 => std_logic_vector(to_unsigned( 16, 8)),5 => std_logic_vector(to_unsigned( 116, 8)),6 => std_logic_vector(to_unsigned( 2, 8)),7 => std_logic_vector(to_unsigned( 7, 8)),8 => std_logic_vector(to_unsigned( 70, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 177) then
				RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),1 => std_logic_vector(to_unsigned( 16, 8)),2 => std_logic_vector(to_unsigned( 50, 8)),3 => std_logic_vector(to_unsigned( 112, 8)),4 => std_logic_vector(to_unsigned( 29, 8)),5 => std_logic_vector(to_unsigned( 61, 8)),6 => std_logic_vector(to_unsigned( 41, 8)),7 => std_logic_vector(to_unsigned( 93, 8)),8 => std_logic_vector(to_unsigned( 107, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 178) then
				RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),1 => std_logic_vector(to_unsigned( 38, 8)),2 => std_logic_vector(to_unsigned( 9, 8)),3 => std_logic_vector(to_unsigned( 92, 8)),4 => std_logic_vector(to_unsigned( 105, 8)),5 => std_logic_vector(to_unsigned( 67, 8)),6 => std_logic_vector(to_unsigned( 22, 8)),7 => std_logic_vector(to_unsigned( 72, 8)),8 => std_logic_vector(to_unsigned( 64, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 179) then
				RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),1 => std_logic_vector(to_unsigned( 11, 8)),2 => std_logic_vector(to_unsigned( 54, 8)),3 => std_logic_vector(to_unsigned( 110, 8)),4 => std_logic_vector(to_unsigned( 69, 8)),5 => std_logic_vector(to_unsigned( 34, 8)),6 => std_logic_vector(to_unsigned( 42, 8)),7 => std_logic_vector(to_unsigned( 58, 8)),8 => std_logic_vector(to_unsigned( 47, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 180) then
				RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),1 => std_logic_vector(to_unsigned( 4, 8)),2 => std_logic_vector(to_unsigned( 120, 8)),3 => std_logic_vector(to_unsigned( 40, 8)),4 => std_logic_vector(to_unsigned( 36, 8)),5 => std_logic_vector(to_unsigned( 114, 8)),6 => std_logic_vector(to_unsigned( 76, 8)),7 => std_logic_vector(to_unsigned( 86, 8)),8 => std_logic_vector(to_unsigned( 84, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 181) then
				RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),1 => std_logic_vector(to_unsigned( 48, 8)),2 => std_logic_vector(to_unsigned( 9, 8)),3 => std_logic_vector(to_unsigned( 22, 8)),4 => std_logic_vector(to_unsigned( 119, 8)),5 => std_logic_vector(to_unsigned( 58, 8)),6 => std_logic_vector(to_unsigned( 115, 8)),7 => std_logic_vector(to_unsigned( 123, 8)),8 => std_logic_vector(to_unsigned( 48, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 182) then
				RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),1 => std_logic_vector(to_unsigned( 49, 8)),2 => std_logic_vector(to_unsigned( 33, 8)),3 => std_logic_vector(to_unsigned( 106, 8)),4 => std_logic_vector(to_unsigned( 54, 8)),5 => std_logic_vector(to_unsigned( 6, 8)),6 => std_logic_vector(to_unsigned( 91, 8)),7 => std_logic_vector(to_unsigned( 25, 8)),8 => std_logic_vector(to_unsigned( 10, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 183) then
				RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),1 => std_logic_vector(to_unsigned( 78, 8)),2 => std_logic_vector(to_unsigned( 26, 8)),3 => std_logic_vector(to_unsigned( 59, 8)),4 => std_logic_vector(to_unsigned( 63, 8)),5 => std_logic_vector(to_unsigned( 36, 8)),6 => std_logic_vector(to_unsigned( 115, 8)),7 => std_logic_vector(to_unsigned( 8, 8)),8 => std_logic_vector(to_unsigned( 92, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 184) then
				RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),1 => std_logic_vector(to_unsigned( 73, 8)),2 => std_logic_vector(to_unsigned( 57, 8)),3 => std_logic_vector(to_unsigned( 87, 8)),4 => std_logic_vector(to_unsigned( 30, 8)),5 => std_logic_vector(to_unsigned( 119, 8)),6 => std_logic_vector(to_unsigned( 68, 8)),7 => std_logic_vector(to_unsigned( 2, 8)),8 => std_logic_vector(to_unsigned( 101, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 185) then
				RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),1 => std_logic_vector(to_unsigned( 91, 8)),2 => std_logic_vector(to_unsigned( 58, 8)),3 => std_logic_vector(to_unsigned( 49, 8)),4 => std_logic_vector(to_unsigned( 75, 8)),5 => std_logic_vector(to_unsigned( 106, 8)),6 => std_logic_vector(to_unsigned( 79, 8)),7 => std_logic_vector(to_unsigned( 18, 8)),8 => std_logic_vector(to_unsigned( 66, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 186) then
				RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),1 => std_logic_vector(to_unsigned( 68, 8)),2 => std_logic_vector(to_unsigned( 122, 8)),3 => std_logic_vector(to_unsigned( 32, 8)),4 => std_logic_vector(to_unsigned( 62, 8)),5 => std_logic_vector(to_unsigned( 12, 8)),6 => std_logic_vector(to_unsigned( 53, 8)),7 => std_logic_vector(to_unsigned( 44, 8)),8 => std_logic_vector(to_unsigned( 113, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 187) then
				RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),1 => std_logic_vector(to_unsigned( 12, 8)),2 => std_logic_vector(to_unsigned( 87, 8)),3 => std_logic_vector(to_unsigned( 19, 8)),4 => std_logic_vector(to_unsigned( 35, 8)),5 => std_logic_vector(to_unsigned( 0, 8)),6 => std_logic_vector(to_unsigned( 80, 8)),7 => std_logic_vector(to_unsigned( 100, 8)),8 => std_logic_vector(to_unsigned( 26, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 188) then
				RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),1 => std_logic_vector(to_unsigned( 49, 8)),2 => std_logic_vector(to_unsigned( 28, 8)),3 => std_logic_vector(to_unsigned( 89, 8)),4 => std_logic_vector(to_unsigned( 43, 8)),5 => std_logic_vector(to_unsigned( 2, 8)),6 => std_logic_vector(to_unsigned( 9, 8)),7 => std_logic_vector(to_unsigned( 63, 8)),8 => std_logic_vector(to_unsigned( 118, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 189) then
				RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),1 => std_logic_vector(to_unsigned( 67, 8)),2 => std_logic_vector(to_unsigned( 83, 8)),3 => std_logic_vector(to_unsigned( 18, 8)),4 => std_logic_vector(to_unsigned( 35, 8)),5 => std_logic_vector(to_unsigned( 93, 8)),6 => std_logic_vector(to_unsigned( 74, 8)),7 => std_logic_vector(to_unsigned( 112, 8)),8 => std_logic_vector(to_unsigned( 87, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 190) then
				RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),1 => std_logic_vector(to_unsigned( 87, 8)),2 => std_logic_vector(to_unsigned( 54, 8)),3 => std_logic_vector(to_unsigned( 61, 8)),4 => std_logic_vector(to_unsigned( 27, 8)),5 => std_logic_vector(to_unsigned( 3, 8)),6 => std_logic_vector(to_unsigned( 116, 8)),7 => std_logic_vector(to_unsigned( 31, 8)),8 => std_logic_vector(to_unsigned( 67, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 191) then
				RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),1 => std_logic_vector(to_unsigned( 40, 8)),2 => std_logic_vector(to_unsigned( 115, 8)),3 => std_logic_vector(to_unsigned( 3, 8)),4 => std_logic_vector(to_unsigned( 26, 8)),5 => std_logic_vector(to_unsigned( 31, 8)),6 => std_logic_vector(to_unsigned( 106, 8)),7 => std_logic_vector(to_unsigned( 76, 8)),8 => std_logic_vector(to_unsigned( 40, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 192) then
				RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),1 => std_logic_vector(to_unsigned( 121, 8)),2 => std_logic_vector(to_unsigned( 75, 8)),3 => std_logic_vector(to_unsigned( 62, 8)),4 => std_logic_vector(to_unsigned( 85, 8)),5 => std_logic_vector(to_unsigned( 81, 8)),6 => std_logic_vector(to_unsigned( 102, 8)),7 => std_logic_vector(to_unsigned( 71, 8)),8 => std_logic_vector(to_unsigned( 108, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 193) then
				RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),1 => std_logic_vector(to_unsigned( 44, 8)),2 => std_logic_vector(to_unsigned( 124, 8)),3 => std_logic_vector(to_unsigned( 21, 8)),4 => std_logic_vector(to_unsigned( 105, 8)),5 => std_logic_vector(to_unsigned( 33, 8)),6 => std_logic_vector(to_unsigned( 9, 8)),7 => std_logic_vector(to_unsigned( 57, 8)),8 => std_logic_vector(to_unsigned( 46, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 194) then
				RAM <= (0 => std_logic_vector(to_unsigned( 115, 8)),1 => std_logic_vector(to_unsigned( 94, 8)),2 => std_logic_vector(to_unsigned( 106, 8)),3 => std_logic_vector(to_unsigned( 35, 8)),4 => std_logic_vector(to_unsigned( 1, 8)),5 => std_logic_vector(to_unsigned( 101, 8)),6 => std_logic_vector(to_unsigned( 21, 8)),7 => std_logic_vector(to_unsigned( 42, 8)),8 => std_logic_vector(to_unsigned( 120, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 195) then
				RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),1 => std_logic_vector(to_unsigned( 46, 8)),2 => std_logic_vector(to_unsigned( 71, 8)),3 => std_logic_vector(to_unsigned( 17, 8)),4 => std_logic_vector(to_unsigned( 26, 8)),5 => std_logic_vector(to_unsigned( 112, 8)),6 => std_logic_vector(to_unsigned( 41, 8)),7 => std_logic_vector(to_unsigned( 82, 8)),8 => std_logic_vector(to_unsigned( 106, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 196) then
				RAM <= (0 => std_logic_vector(to_unsigned( 28, 8)),1 => std_logic_vector(to_unsigned( 64, 8)),2 => std_logic_vector(to_unsigned( 78, 8)),3 => std_logic_vector(to_unsigned( 53, 8)),4 => std_logic_vector(to_unsigned( 37, 8)),5 => std_logic_vector(to_unsigned( 6, 8)),6 => std_logic_vector(to_unsigned( 16, 8)),7 => std_logic_vector(to_unsigned( 82, 8)),8 => std_logic_vector(to_unsigned( 76, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 197) then
				RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),1 => std_logic_vector(to_unsigned( 35, 8)),2 => std_logic_vector(to_unsigned( 31, 8)),3 => std_logic_vector(to_unsigned( 87, 8)),4 => std_logic_vector(to_unsigned( 97, 8)),5 => std_logic_vector(to_unsigned( 106, 8)),6 => std_logic_vector(to_unsigned( 118, 8)),7 => std_logic_vector(to_unsigned( 22, 8)),8 => std_logic_vector(to_unsigned( 4, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 198) then
				RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),1 => std_logic_vector(to_unsigned( 92, 8)),2 => std_logic_vector(to_unsigned( 75, 8)),3 => std_logic_vector(to_unsigned( 30, 8)),4 => std_logic_vector(to_unsigned( 66, 8)),5 => std_logic_vector(to_unsigned( 16, 8)),6 => std_logic_vector(to_unsigned( 52, 8)),7 => std_logic_vector(to_unsigned( 109, 8)),8 => std_logic_vector(to_unsigned( 20, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 199) then
				RAM <= (0 => std_logic_vector(to_unsigned( 90, 8)),1 => std_logic_vector(to_unsigned( 10, 8)),2 => std_logic_vector(to_unsigned( 30, 8)),3 => std_logic_vector(to_unsigned( 0, 8)),4 => std_logic_vector(to_unsigned( 46, 8)),5 => std_logic_vector(to_unsigned( 77, 8)),6 => std_logic_vector(to_unsigned( 70, 8)),7 => std_logic_vector(to_unsigned( 54, 8)),8 => std_logic_vector(to_unsigned( 107, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 200) then
				RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),1 => std_logic_vector(to_unsigned( 59, 8)),2 => std_logic_vector(to_unsigned( 48, 8)),3 => std_logic_vector(to_unsigned( 75, 8)),4 => std_logic_vector(to_unsigned( 104, 8)),5 => std_logic_vector(to_unsigned( 38, 8)),6 => std_logic_vector(to_unsigned( 111, 8)),7 => std_logic_vector(to_unsigned( 64, 8)),8 => std_logic_vector(to_unsigned( 58, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 201) then
				RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),1 => std_logic_vector(to_unsigned( 34, 8)),2 => std_logic_vector(to_unsigned( 97, 8)),3 => std_logic_vector(to_unsigned( 56, 8)),4 => std_logic_vector(to_unsigned( 115, 8)),5 => std_logic_vector(to_unsigned( 0, 8)),6 => std_logic_vector(to_unsigned( 82, 8)),7 => std_logic_vector(to_unsigned( 4, 8)),8 => std_logic_vector(to_unsigned( 101, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 202) then
				RAM <= (0 => std_logic_vector(to_unsigned( 86, 8)),1 => std_logic_vector(to_unsigned( 33, 8)),2 => std_logic_vector(to_unsigned( 10, 8)),3 => std_logic_vector(to_unsigned( 62, 8)),4 => std_logic_vector(to_unsigned( 24, 8)),5 => std_logic_vector(to_unsigned( 19, 8)),6 => std_logic_vector(to_unsigned( 96, 8)),7 => std_logic_vector(to_unsigned( 109, 8)),8 => std_logic_vector(to_unsigned( 116, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 203) then
				RAM <= (0 => std_logic_vector(to_unsigned( 77, 8)),1 => std_logic_vector(to_unsigned( 21, 8)),2 => std_logic_vector(to_unsigned( 27, 8)),3 => std_logic_vector(to_unsigned( 109, 8)),4 => std_logic_vector(to_unsigned( 60, 8)),5 => std_logic_vector(to_unsigned( 8, 8)),6 => std_logic_vector(to_unsigned( 40, 8)),7 => std_logic_vector(to_unsigned( 82, 8)),8 => std_logic_vector(to_unsigned( 77, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 204) then
				RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),1 => std_logic_vector(to_unsigned( 74, 8)),2 => std_logic_vector(to_unsigned( 38, 8)),3 => std_logic_vector(to_unsigned( 99, 8)),4 => std_logic_vector(to_unsigned( 25, 8)),5 => std_logic_vector(to_unsigned( 20, 8)),6 => std_logic_vector(to_unsigned( 70, 8)),7 => std_logic_vector(to_unsigned( 86, 8)),8 => std_logic_vector(to_unsigned( 22, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 205) then
				RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),1 => std_logic_vector(to_unsigned( 47, 8)),2 => std_logic_vector(to_unsigned( 79, 8)),3 => std_logic_vector(to_unsigned( 23, 8)),4 => std_logic_vector(to_unsigned( 75, 8)),5 => std_logic_vector(to_unsigned( 37, 8)),6 => std_logic_vector(to_unsigned( 108, 8)),7 => std_logic_vector(to_unsigned( 41, 8)),8 => std_logic_vector(to_unsigned( 31, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 206) then
				RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),1 => std_logic_vector(to_unsigned( 104, 8)),2 => std_logic_vector(to_unsigned( 12, 8)),3 => std_logic_vector(to_unsigned( 123, 8)),4 => std_logic_vector(to_unsigned( 67, 8)),5 => std_logic_vector(to_unsigned( 111, 8)),6 => std_logic_vector(to_unsigned( 88, 8)),7 => std_logic_vector(to_unsigned( 60, 8)),8 => std_logic_vector(to_unsigned( 70, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 207) then
				RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),1 => std_logic_vector(to_unsigned( 52, 8)),2 => std_logic_vector(to_unsigned( 67, 8)),3 => std_logic_vector(to_unsigned( 118, 8)),4 => std_logic_vector(to_unsigned( 124, 8)),5 => std_logic_vector(to_unsigned( 112, 8)),6 => std_logic_vector(to_unsigned( 33, 8)),7 => std_logic_vector(to_unsigned( 81, 8)),8 => std_logic_vector(to_unsigned( 117, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 208) then
				RAM <= (0 => std_logic_vector(to_unsigned( 56, 8)),1 => std_logic_vector(to_unsigned( 118, 8)),2 => std_logic_vector(to_unsigned( 28, 8)),3 => std_logic_vector(to_unsigned( 40, 8)),4 => std_logic_vector(to_unsigned( 67, 8)),5 => std_logic_vector(to_unsigned( 24, 8)),6 => std_logic_vector(to_unsigned( 92, 8)),7 => std_logic_vector(to_unsigned( 102, 8)),8 => std_logic_vector(to_unsigned( 34, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 209) then
				RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),1 => std_logic_vector(to_unsigned( 40, 8)),2 => std_logic_vector(to_unsigned( 48, 8)),3 => std_logic_vector(to_unsigned( 34, 8)),4 => std_logic_vector(to_unsigned( 88, 8)),5 => std_logic_vector(to_unsigned( 97, 8)),6 => std_logic_vector(to_unsigned( 101, 8)),7 => std_logic_vector(to_unsigned( 121, 8)),8 => std_logic_vector(to_unsigned( 28, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 210) then
				RAM <= (0 => std_logic_vector(to_unsigned( 87, 8)),1 => std_logic_vector(to_unsigned( 112, 8)),2 => std_logic_vector(to_unsigned( 16, 8)),3 => std_logic_vector(to_unsigned( 68, 8)),4 => std_logic_vector(to_unsigned( 52, 8)),5 => std_logic_vector(to_unsigned( 43, 8)),6 => std_logic_vector(to_unsigned( 72, 8)),7 => std_logic_vector(to_unsigned( 91, 8)),8 => std_logic_vector(to_unsigned( 98, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 211) then
				RAM <= (0 => std_logic_vector(to_unsigned( 15, 8)),1 => std_logic_vector(to_unsigned( 58, 8)),2 => std_logic_vector(to_unsigned( 38, 8)),3 => std_logic_vector(to_unsigned( 106, 8)),4 => std_logic_vector(to_unsigned( 62, 8)),5 => std_logic_vector(to_unsigned( 25, 8)),6 => std_logic_vector(to_unsigned( 42, 8)),7 => std_logic_vector(to_unsigned( 66, 8)),8 => std_logic_vector(to_unsigned( 6, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 212) then
				RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),1 => std_logic_vector(to_unsigned( 20, 8)),2 => std_logic_vector(to_unsigned( 103, 8)),3 => std_logic_vector(to_unsigned( 122, 8)),4 => std_logic_vector(to_unsigned( 39, 8)),5 => std_logic_vector(to_unsigned( 84, 8)),6 => std_logic_vector(to_unsigned( 34, 8)),7 => std_logic_vector(to_unsigned( 50, 8)),8 => std_logic_vector(to_unsigned( 60, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 213) then
				RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),1 => std_logic_vector(to_unsigned( 81, 8)),2 => std_logic_vector(to_unsigned( 124, 8)),3 => std_logic_vector(to_unsigned( 104, 8)),4 => std_logic_vector(to_unsigned( 75, 8)),5 => std_logic_vector(to_unsigned( 10, 8)),6 => std_logic_vector(to_unsigned( 85, 8)),7 => std_logic_vector(to_unsigned( 45, 8)),8 => std_logic_vector(to_unsigned( 124, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 214) then
				RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),1 => std_logic_vector(to_unsigned( 57, 8)),2 => std_logic_vector(to_unsigned( 27, 8)),3 => std_logic_vector(to_unsigned( 8, 8)),4 => std_logic_vector(to_unsigned( 16, 8)),5 => std_logic_vector(to_unsigned( 89, 8)),6 => std_logic_vector(to_unsigned( 111, 8)),7 => std_logic_vector(to_unsigned( 124, 8)),8 => std_logic_vector(to_unsigned( 22, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 215) then
				RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),1 => std_logic_vector(to_unsigned( 88, 8)),2 => std_logic_vector(to_unsigned( 12, 8)),3 => std_logic_vector(to_unsigned( 113, 8)),4 => std_logic_vector(to_unsigned( 17, 8)),5 => std_logic_vector(to_unsigned( 54, 8)),6 => std_logic_vector(to_unsigned( 26, 8)),7 => std_logic_vector(to_unsigned( 98, 8)),8 => std_logic_vector(to_unsigned( 57, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 216) then
				RAM <= (0 => std_logic_vector(to_unsigned( 47, 8)),1 => std_logic_vector(to_unsigned( 34, 8)),2 => std_logic_vector(to_unsigned( 109, 8)),3 => std_logic_vector(to_unsigned( 101, 8)),4 => std_logic_vector(to_unsigned( 21, 8)),5 => std_logic_vector(to_unsigned( 54, 8)),6 => std_logic_vector(to_unsigned( 116, 8)),7 => std_logic_vector(to_unsigned( 87, 8)),8 => std_logic_vector(to_unsigned( 28, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 217) then
				RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),1 => std_logic_vector(to_unsigned( 12, 8)),2 => std_logic_vector(to_unsigned( 44, 8)),3 => std_logic_vector(to_unsigned( 6, 8)),4 => std_logic_vector(to_unsigned( 18, 8)),5 => std_logic_vector(to_unsigned( 27, 8)),6 => std_logic_vector(to_unsigned( 115, 8)),7 => std_logic_vector(to_unsigned( 75, 8)),8 => std_logic_vector(to_unsigned( 49, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 218) then
				RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),1 => std_logic_vector(to_unsigned( 36, 8)),2 => std_logic_vector(to_unsigned( 85, 8)),3 => std_logic_vector(to_unsigned( 95, 8)),4 => std_logic_vector(to_unsigned( 5, 8)),5 => std_logic_vector(to_unsigned( 69, 8)),6 => std_logic_vector(to_unsigned( 75, 8)),7 => std_logic_vector(to_unsigned( 16, 8)),8 => std_logic_vector(to_unsigned( 69, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 219) then
				RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),1 => std_logic_vector(to_unsigned( 60, 8)),2 => std_logic_vector(to_unsigned( 4, 8)),3 => std_logic_vector(to_unsigned( 77, 8)),4 => std_logic_vector(to_unsigned( 34, 8)),5 => std_logic_vector(to_unsigned( 110, 8)),6 => std_logic_vector(to_unsigned( 23, 8)),7 => std_logic_vector(to_unsigned( 54, 8)),8 => std_logic_vector(to_unsigned( 27, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 220) then
				RAM <= (0 => std_logic_vector(to_unsigned( 70, 8)),1 => std_logic_vector(to_unsigned( 21, 8)),2 => std_logic_vector(to_unsigned( 39, 8)),3 => std_logic_vector(to_unsigned( 120, 8)),4 => std_logic_vector(to_unsigned( 102, 8)),5 => std_logic_vector(to_unsigned( 87, 8)),6 => std_logic_vector(to_unsigned( 0, 8)),7 => std_logic_vector(to_unsigned( 11, 8)),8 => std_logic_vector(to_unsigned( 43, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 221) then
				RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),1 => std_logic_vector(to_unsigned( 87, 8)),2 => std_logic_vector(to_unsigned( 47, 8)),3 => std_logic_vector(to_unsigned( 109, 8)),4 => std_logic_vector(to_unsigned( 75, 8)),5 => std_logic_vector(to_unsigned( 61, 8)),6 => std_logic_vector(to_unsigned( 41, 8)),7 => std_logic_vector(to_unsigned( 56, 8)),8 => std_logic_vector(to_unsigned( 110, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 222) then
				RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),1 => std_logic_vector(to_unsigned( 30, 8)),2 => std_logic_vector(to_unsigned( 14, 8)),3 => std_logic_vector(to_unsigned( 46, 8)),4 => std_logic_vector(to_unsigned( 60, 8)),5 => std_logic_vector(to_unsigned( 5, 8)),6 => std_logic_vector(to_unsigned( 78, 8)),7 => std_logic_vector(to_unsigned( 105, 8)),8 => std_logic_vector(to_unsigned( 74, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 223) then
				RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),1 => std_logic_vector(to_unsigned( 7, 8)),2 => std_logic_vector(to_unsigned( 69, 8)),3 => std_logic_vector(to_unsigned( 48, 8)),4 => std_logic_vector(to_unsigned( 115, 8)),5 => std_logic_vector(to_unsigned( 101, 8)),6 => std_logic_vector(to_unsigned( 42, 8)),7 => std_logic_vector(to_unsigned( 75, 8)),8 => std_logic_vector(to_unsigned( 106, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 224) then
				RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),1 => std_logic_vector(to_unsigned( 3, 8)),2 => std_logic_vector(to_unsigned( 94, 8)),3 => std_logic_vector(to_unsigned( 77, 8)),4 => std_logic_vector(to_unsigned( 59, 8)),5 => std_logic_vector(to_unsigned( 83, 8)),6 => std_logic_vector(to_unsigned( 20, 8)),7 => std_logic_vector(to_unsigned( 49, 8)),8 => std_logic_vector(to_unsigned( 25, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 225) then
				RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),1 => std_logic_vector(to_unsigned( 60, 8)),2 => std_logic_vector(to_unsigned( 81, 8)),3 => std_logic_vector(to_unsigned( 69, 8)),4 => std_logic_vector(to_unsigned( 96, 8)),5 => std_logic_vector(to_unsigned( 9, 8)),6 => std_logic_vector(to_unsigned( 26, 8)),7 => std_logic_vector(to_unsigned( 88, 8)),8 => std_logic_vector(to_unsigned( 118, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 226) then
				RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),1 => std_logic_vector(to_unsigned( 17, 8)),2 => std_logic_vector(to_unsigned( 38, 8)),3 => std_logic_vector(to_unsigned( 71, 8)),4 => std_logic_vector(to_unsigned( 113, 8)),5 => std_logic_vector(to_unsigned( 60, 8)),6 => std_logic_vector(to_unsigned( 8, 8)),7 => std_logic_vector(to_unsigned( 120, 8)),8 => std_logic_vector(to_unsigned( 127, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 227) then
				RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),1 => std_logic_vector(to_unsigned( 118, 8)),2 => std_logic_vector(to_unsigned( 4, 8)),3 => std_logic_vector(to_unsigned( 40, 8)),4 => std_logic_vector(to_unsigned( 107, 8)),5 => std_logic_vector(to_unsigned( 101, 8)),6 => std_logic_vector(to_unsigned( 20, 8)),7 => std_logic_vector(to_unsigned( 36, 8)),8 => std_logic_vector(to_unsigned( 33, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 228) then
				RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),1 => std_logic_vector(to_unsigned( 54, 8)),2 => std_logic_vector(to_unsigned( 45, 8)),3 => std_logic_vector(to_unsigned( 12, 8)),4 => std_logic_vector(to_unsigned( 86, 8)),5 => std_logic_vector(to_unsigned( 76, 8)),6 => std_logic_vector(to_unsigned( 72, 8)),7 => std_logic_vector(to_unsigned( 37, 8)),8 => std_logic_vector(to_unsigned( 0, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 229) then
				RAM <= (0 => std_logic_vector(to_unsigned( 91, 8)),1 => std_logic_vector(to_unsigned( 108, 8)),2 => std_logic_vector(to_unsigned( 87, 8)),3 => std_logic_vector(to_unsigned( 0, 8)),4 => std_logic_vector(to_unsigned( 42, 8)),5 => std_logic_vector(to_unsigned( 81, 8)),6 => std_logic_vector(to_unsigned( 26, 8)),7 => std_logic_vector(to_unsigned( 47, 8)),8 => std_logic_vector(to_unsigned( 93, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 230) then
				RAM <= (0 => std_logic_vector(to_unsigned( 27, 8)),1 => std_logic_vector(to_unsigned( 12, 8)),2 => std_logic_vector(to_unsigned( 21, 8)),3 => std_logic_vector(to_unsigned( 99, 8)),4 => std_logic_vector(to_unsigned( 106, 8)),5 => std_logic_vector(to_unsigned( 67, 8)),6 => std_logic_vector(to_unsigned( 92, 8)),7 => std_logic_vector(to_unsigned( 4, 8)),8 => std_logic_vector(to_unsigned( 20, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 231) then
				RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),1 => std_logic_vector(to_unsigned( 94, 8)),2 => std_logic_vector(to_unsigned( 40, 8)),3 => std_logic_vector(to_unsigned( 12, 8)),4 => std_logic_vector(to_unsigned( 2, 8)),5 => std_logic_vector(to_unsigned( 118, 8)),6 => std_logic_vector(to_unsigned( 71, 8)),7 => std_logic_vector(to_unsigned( 33, 8)),8 => std_logic_vector(to_unsigned( 7, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 232) then
				RAM <= (0 => std_logic_vector(to_unsigned( 109, 8)),1 => std_logic_vector(to_unsigned( 6, 8)),2 => std_logic_vector(to_unsigned( 43, 8)),3 => std_logic_vector(to_unsigned( 104, 8)),4 => std_logic_vector(to_unsigned( 87, 8)),5 => std_logic_vector(to_unsigned( 118, 8)),6 => std_logic_vector(to_unsigned( 114, 8)),7 => std_logic_vector(to_unsigned( 60, 8)),8 => std_logic_vector(to_unsigned( 5, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 233) then
				RAM <= (0 => std_logic_vector(to_unsigned( 41, 8)),1 => std_logic_vector(to_unsigned( 55, 8)),2 => std_logic_vector(to_unsigned( 29, 8)),3 => std_logic_vector(to_unsigned( 77, 8)),4 => std_logic_vector(to_unsigned( 90, 8)),5 => std_logic_vector(to_unsigned( 116, 8)),6 => std_logic_vector(to_unsigned( 70, 8)),7 => std_logic_vector(to_unsigned( 86, 8)),8 => std_logic_vector(to_unsigned( 55, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 234) then
				RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),1 => std_logic_vector(to_unsigned( 84, 8)),2 => std_logic_vector(to_unsigned( 60, 8)),3 => std_logic_vector(to_unsigned( 96, 8)),4 => std_logic_vector(to_unsigned( 23, 8)),5 => std_logic_vector(to_unsigned( 47, 8)),6 => std_logic_vector(to_unsigned( 103, 8)),7 => std_logic_vector(to_unsigned( 39, 8)),8 => std_logic_vector(to_unsigned( 43, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 235) then
				RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),1 => std_logic_vector(to_unsigned( 21, 8)),2 => std_logic_vector(to_unsigned( 9, 8)),3 => std_logic_vector(to_unsigned( 3, 8)),4 => std_logic_vector(to_unsigned( 121, 8)),5 => std_logic_vector(to_unsigned( 98, 8)),6 => std_logic_vector(to_unsigned( 92, 8)),7 => std_logic_vector(to_unsigned( 70, 8)),8 => std_logic_vector(to_unsigned( 3, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 236) then
				RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),1 => std_logic_vector(to_unsigned( 122, 8)),2 => std_logic_vector(to_unsigned( 31, 8)),3 => std_logic_vector(to_unsigned( 49, 8)),4 => std_logic_vector(to_unsigned( 101, 8)),5 => std_logic_vector(to_unsigned( 117, 8)),6 => std_logic_vector(to_unsigned( 13, 8)),7 => std_logic_vector(to_unsigned( 72, 8)),8 => std_logic_vector(to_unsigned( 122, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 237) then
				RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),1 => std_logic_vector(to_unsigned( 43, 8)),2 => std_logic_vector(to_unsigned( 59, 8)),3 => std_logic_vector(to_unsigned( 76, 8)),4 => std_logic_vector(to_unsigned( 17, 8)),5 => std_logic_vector(to_unsigned( 26, 8)),6 => std_logic_vector(to_unsigned( 65, 8)),7 => std_logic_vector(to_unsigned( 96, 8)),8 => std_logic_vector(to_unsigned( 89, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 238) then
				RAM <= (0 => std_logic_vector(to_unsigned( 29, 8)),1 => std_logic_vector(to_unsigned( 83, 8)),2 => std_logic_vector(to_unsigned( 105, 8)),3 => std_logic_vector(to_unsigned( 47, 8)),4 => std_logic_vector(to_unsigned( 23, 8)),5 => std_logic_vector(to_unsigned( 60, 8)),6 => std_logic_vector(to_unsigned( 72, 8)),7 => std_logic_vector(to_unsigned( 124, 8)),8 => std_logic_vector(to_unsigned( 63, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 239) then
				RAM <= (0 => std_logic_vector(to_unsigned( 112, 8)),1 => std_logic_vector(to_unsigned( 65, 8)),2 => std_logic_vector(to_unsigned( 99, 8)),3 => std_logic_vector(to_unsigned( 38, 8)),4 => std_logic_vector(to_unsigned( 51, 8)),5 => std_logic_vector(to_unsigned( 3, 8)),6 => std_logic_vector(to_unsigned( 94, 8)),7 => std_logic_vector(to_unsigned( 108, 8)),8 => std_logic_vector(to_unsigned( 111, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 240) then
				RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),1 => std_logic_vector(to_unsigned( 30, 8)),2 => std_logic_vector(to_unsigned( 24, 8)),3 => std_logic_vector(to_unsigned( 113, 8)),4 => std_logic_vector(to_unsigned( 58, 8)),5 => std_logic_vector(to_unsigned( 7, 8)),6 => std_logic_vector(to_unsigned( 66, 8)),7 => std_logic_vector(to_unsigned( 102, 8)),8 => std_logic_vector(to_unsigned( 95, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 241) then
				RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),1 => std_logic_vector(to_unsigned( 100, 8)),2 => std_logic_vector(to_unsigned( 25, 8)),3 => std_logic_vector(to_unsigned( 36, 8)),4 => std_logic_vector(to_unsigned( 2, 8)),5 => std_logic_vector(to_unsigned( 85, 8)),6 => std_logic_vector(to_unsigned( 64, 8)),7 => std_logic_vector(to_unsigned( 124, 8)),8 => std_logic_vector(to_unsigned( 13, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 242) then
				RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),1 => std_logic_vector(to_unsigned( 70, 8)),2 => std_logic_vector(to_unsigned( 62, 8)),3 => std_logic_vector(to_unsigned( 119, 8)),4 => std_logic_vector(to_unsigned( 41, 8)),5 => std_logic_vector(to_unsigned( 108, 8)),6 => std_logic_vector(to_unsigned( 95, 8)),7 => std_logic_vector(to_unsigned( 49, 8)),8 => std_logic_vector(to_unsigned( 79, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 243) then
				RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),1 => std_logic_vector(to_unsigned( 94, 8)),2 => std_logic_vector(to_unsigned( 75, 8)),3 => std_logic_vector(to_unsigned( 87, 8)),4 => std_logic_vector(to_unsigned( 111, 8)),5 => std_logic_vector(to_unsigned( 116, 8)),6 => std_logic_vector(to_unsigned( 63, 8)),7 => std_logic_vector(to_unsigned( 26, 8)),8 => std_logic_vector(to_unsigned( 12, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 244) then
				RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),1 => std_logic_vector(to_unsigned( 123, 8)),2 => std_logic_vector(to_unsigned( 75, 8)),3 => std_logic_vector(to_unsigned( 47, 8)),4 => std_logic_vector(to_unsigned( 14, 8)),5 => std_logic_vector(to_unsigned( 119, 8)),6 => std_logic_vector(to_unsigned( 59, 8)),7 => std_logic_vector(to_unsigned( 23, 8)),8 => std_logic_vector(to_unsigned( 64, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 245) then
				RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),1 => std_logic_vector(to_unsigned( 103, 8)),2 => std_logic_vector(to_unsigned( 2, 8)),3 => std_logic_vector(to_unsigned( 123, 8)),4 => std_logic_vector(to_unsigned( 44, 8)),5 => std_logic_vector(to_unsigned( 118, 8)),6 => std_logic_vector(to_unsigned( 97, 8)),7 => std_logic_vector(to_unsigned( 16, 8)),8 => std_logic_vector(to_unsigned( 48, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 246) then
				RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),1 => std_logic_vector(to_unsigned( 1, 8)),2 => std_logic_vector(to_unsigned( 24, 8)),3 => std_logic_vector(to_unsigned( 44, 8)),4 => std_logic_vector(to_unsigned( 37, 8)),5 => std_logic_vector(to_unsigned( 13, 8)),6 => std_logic_vector(to_unsigned( 83, 8)),7 => std_logic_vector(to_unsigned( 60, 8)),8 => std_logic_vector(to_unsigned( 98, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 247) then
				RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),1 => std_logic_vector(to_unsigned( 80, 8)),2 => std_logic_vector(to_unsigned( 124, 8)),3 => std_logic_vector(to_unsigned( 48, 8)),4 => std_logic_vector(to_unsigned( 71, 8)),5 => std_logic_vector(to_unsigned( 62, 8)),6 => std_logic_vector(to_unsigned( 43, 8)),7 => std_logic_vector(to_unsigned( 0, 8)),8 => std_logic_vector(to_unsigned( 52, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 248) then
				RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),1 => std_logic_vector(to_unsigned( 58, 8)),2 => std_logic_vector(to_unsigned( 39, 8)),3 => std_logic_vector(to_unsigned( 105, 8)),4 => std_logic_vector(to_unsigned( 123, 8)),5 => std_logic_vector(to_unsigned( 30, 8)),6 => std_logic_vector(to_unsigned( 12, 8)),7 => std_logic_vector(to_unsigned( 92, 8)),8 => std_logic_vector(to_unsigned( 77, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 249) then
				RAM <= (0 => std_logic_vector(to_unsigned( 53, 8)),1 => std_logic_vector(to_unsigned( 60, 8)),2 => std_logic_vector(to_unsigned( 9, 8)),3 => std_logic_vector(to_unsigned( 73, 8)),4 => std_logic_vector(to_unsigned( 92, 8)),5 => std_logic_vector(to_unsigned( 13, 8)),6 => std_logic_vector(to_unsigned( 1, 8)),7 => std_logic_vector(to_unsigned( 26, 8)),8 => std_logic_vector(to_unsigned( 52, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 250) then
				RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),1 => std_logic_vector(to_unsigned( 11, 8)),2 => std_logic_vector(to_unsigned( 64, 8)),3 => std_logic_vector(to_unsigned( 109, 8)),4 => std_logic_vector(to_unsigned( 92, 8)),5 => std_logic_vector(to_unsigned( 69, 8)),6 => std_logic_vector(to_unsigned( 50, 8)),7 => std_logic_vector(to_unsigned( 44, 8)),8 => std_logic_vector(to_unsigned( 59, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 251) then
				RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),1 => std_logic_vector(to_unsigned( 73, 8)),2 => std_logic_vector(to_unsigned( 34, 8)),3 => std_logic_vector(to_unsigned( 5, 8)),4 => std_logic_vector(to_unsigned( 63, 8)),5 => std_logic_vector(to_unsigned( 117, 8)),6 => std_logic_vector(to_unsigned( 20, 8)),7 => std_logic_vector(to_unsigned( 107, 8)),8 => std_logic_vector(to_unsigned( 77, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 252) then
				RAM <= (0 => std_logic_vector(to_unsigned( 26, 8)),1 => std_logic_vector(to_unsigned( 4, 8)),2 => std_logic_vector(to_unsigned( 37, 8)),3 => std_logic_vector(to_unsigned( 81, 8)),4 => std_logic_vector(to_unsigned( 50, 8)),5 => std_logic_vector(to_unsigned( 41, 8)),6 => std_logic_vector(to_unsigned( 89, 8)),7 => std_logic_vector(to_unsigned( 104, 8)),8 => std_logic_vector(to_unsigned( 112, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 253) then
				RAM <= (0 => std_logic_vector(to_unsigned( 77, 8)),1 => std_logic_vector(to_unsigned( 37, 8)),2 => std_logic_vector(to_unsigned( 57, 8)),3 => std_logic_vector(to_unsigned( 26, 8)),4 => std_logic_vector(to_unsigned( 83, 8)),5 => std_logic_vector(to_unsigned( 95, 8)),6 => std_logic_vector(to_unsigned( 102, 8)),7 => std_logic_vector(to_unsigned( 67, 8)),8 => std_logic_vector(to_unsigned( 52, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 254) then
				RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),1 => std_logic_vector(to_unsigned( 57, 8)),2 => std_logic_vector(to_unsigned( 15, 8)),3 => std_logic_vector(to_unsigned( 105, 8)),4 => std_logic_vector(to_unsigned( 3, 8)),5 => std_logic_vector(to_unsigned( 35, 8)),6 => std_logic_vector(to_unsigned( 86, 8)),7 => std_logic_vector(to_unsigned( 122, 8)),8 => std_logic_vector(to_unsigned( 72, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 255) then
				RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),1 => std_logic_vector(to_unsigned( 30, 8)),2 => std_logic_vector(to_unsigned( 90, 8)),3 => std_logic_vector(to_unsigned( 71, 8)),4 => std_logic_vector(to_unsigned( 16, 8)),5 => std_logic_vector(to_unsigned( 57, 8)),6 => std_logic_vector(to_unsigned( 37, 8)),7 => std_logic_vector(to_unsigned( 62, 8)),8 => std_logic_vector(to_unsigned( 42, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 256) then
				RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),1 => std_logic_vector(to_unsigned( 50, 8)),2 => std_logic_vector(to_unsigned( 55, 8)),3 => std_logic_vector(to_unsigned( 3, 8)),4 => std_logic_vector(to_unsigned( 92, 8)),5 => std_logic_vector(to_unsigned( 11, 8)),6 => std_logic_vector(to_unsigned( 36, 8)),7 => std_logic_vector(to_unsigned( 16, 8)),8 => std_logic_vector(to_unsigned( 80, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 257) then
				RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),1 => std_logic_vector(to_unsigned( 13, 8)),2 => std_logic_vector(to_unsigned( 70, 8)),3 => std_logic_vector(to_unsigned( 75, 8)),4 => std_logic_vector(to_unsigned( 41, 8)),5 => std_logic_vector(to_unsigned( 29, 8)),6 => std_logic_vector(to_unsigned( 123, 8)),7 => std_logic_vector(to_unsigned( 48, 8)),8 => std_logic_vector(to_unsigned( 23, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 258) then
				RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),1 => std_logic_vector(to_unsigned( 19, 8)),2 => std_logic_vector(to_unsigned( 85, 8)),3 => std_logic_vector(to_unsigned( 108, 8)),4 => std_logic_vector(to_unsigned( 62, 8)),5 => std_logic_vector(to_unsigned( 0, 8)),6 => std_logic_vector(to_unsigned( 57, 8)),7 => std_logic_vector(to_unsigned( 100, 8)),8 => std_logic_vector(to_unsigned( 120, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 259) then
				RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),1 => std_logic_vector(to_unsigned( 39, 8)),2 => std_logic_vector(to_unsigned( 108, 8)),3 => std_logic_vector(to_unsigned( 45, 8)),4 => std_logic_vector(to_unsigned( 27, 8)),5 => std_logic_vector(to_unsigned( 87, 8)),6 => std_logic_vector(to_unsigned( 16, 8)),7 => std_logic_vector(to_unsigned( 75, 8)),8 => std_logic_vector(to_unsigned( 3, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 260) then
				RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),1 => std_logic_vector(to_unsigned( 69, 8)),2 => std_logic_vector(to_unsigned( 10, 8)),3 => std_logic_vector(to_unsigned( 35, 8)),4 => std_logic_vector(to_unsigned( 56, 8)),5 => std_logic_vector(to_unsigned( 86, 8)),6 => std_logic_vector(to_unsigned( 2, 8)),7 => std_logic_vector(to_unsigned( 114, 8)),8 => std_logic_vector(to_unsigned( 104, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 261) then
				RAM <= (0 => std_logic_vector(to_unsigned( 114, 8)),1 => std_logic_vector(to_unsigned( 96, 8)),2 => std_logic_vector(to_unsigned( 108, 8)),3 => std_logic_vector(to_unsigned( 54, 8)),4 => std_logic_vector(to_unsigned( 83, 8)),5 => std_logic_vector(to_unsigned( 42, 8)),6 => std_logic_vector(to_unsigned( 9, 8)),7 => std_logic_vector(to_unsigned( 104, 8)),8 => std_logic_vector(to_unsigned( 74, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 262) then
				RAM <= (0 => std_logic_vector(to_unsigned( 92, 8)),1 => std_logic_vector(to_unsigned( 18, 8)),2 => std_logic_vector(to_unsigned( 80, 8)),3 => std_logic_vector(to_unsigned( 29, 8)),4 => std_logic_vector(to_unsigned( 113, 8)),5 => std_logic_vector(to_unsigned( 58, 8)),6 => std_logic_vector(to_unsigned( 11, 8)),7 => std_logic_vector(to_unsigned( 52, 8)),8 => std_logic_vector(to_unsigned( 122, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 263) then
				RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),1 => std_logic_vector(to_unsigned( 104, 8)),2 => std_logic_vector(to_unsigned( 110, 8)),3 => std_logic_vector(to_unsigned( 49, 8)),4 => std_logic_vector(to_unsigned( 15, 8)),5 => std_logic_vector(to_unsigned( 27, 8)),6 => std_logic_vector(to_unsigned( 41, 8)),7 => std_logic_vector(to_unsigned( 72, 8)),8 => std_logic_vector(to_unsigned( 117, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 264) then
				RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),1 => std_logic_vector(to_unsigned( 76, 8)),2 => std_logic_vector(to_unsigned( 65, 8)),3 => std_logic_vector(to_unsigned( 106, 8)),4 => std_logic_vector(to_unsigned( 29, 8)),5 => std_logic_vector(to_unsigned( 23, 8)),6 => std_logic_vector(to_unsigned( 0, 8)),7 => std_logic_vector(to_unsigned( 58, 8)),8 => std_logic_vector(to_unsigned( 29, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 265) then
				RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),1 => std_logic_vector(to_unsigned( 45, 8)),2 => std_logic_vector(to_unsigned( 70, 8)),3 => std_logic_vector(to_unsigned( 6, 8)),4 => std_logic_vector(to_unsigned( 11, 8)),5 => std_logic_vector(to_unsigned( 58, 8)),6 => std_logic_vector(to_unsigned( 24, 8)),7 => std_logic_vector(to_unsigned( 49, 8)),8 => std_logic_vector(to_unsigned( 51, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 266) then
				RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),1 => std_logic_vector(to_unsigned( 122, 8)),2 => std_logic_vector(to_unsigned( 109, 8)),3 => std_logic_vector(to_unsigned( 41, 8)),4 => std_logic_vector(to_unsigned( 69, 8)),5 => std_logic_vector(to_unsigned( 14, 8)),6 => std_logic_vector(to_unsigned( 32, 8)),7 => std_logic_vector(to_unsigned( 22, 8)),8 => std_logic_vector(to_unsigned( 22, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 267) then
				RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),1 => std_logic_vector(to_unsigned( 49, 8)),2 => std_logic_vector(to_unsigned( 101, 8)),3 => std_logic_vector(to_unsigned( 68, 8)),4 => std_logic_vector(to_unsigned( 92, 8)),5 => std_logic_vector(to_unsigned( 76, 8)),6 => std_logic_vector(to_unsigned( 30, 8)),7 => std_logic_vector(to_unsigned( 110, 8)),8 => std_logic_vector(to_unsigned( 98, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 268) then
				RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),1 => std_logic_vector(to_unsigned( 65, 8)),2 => std_logic_vector(to_unsigned( 90, 8)),3 => std_logic_vector(to_unsigned( 121, 8)),4 => std_logic_vector(to_unsigned( 29, 8)),5 => std_logic_vector(to_unsigned( 54, 8)),6 => std_logic_vector(to_unsigned( 78, 8)),7 => std_logic_vector(to_unsigned( 85, 8)),8 => std_logic_vector(to_unsigned( 97, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 269) then
				RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),1 => std_logic_vector(to_unsigned( 121, 8)),2 => std_logic_vector(to_unsigned( 14, 8)),3 => std_logic_vector(to_unsigned( 61, 8)),4 => std_logic_vector(to_unsigned( 96, 8)),5 => std_logic_vector(to_unsigned( 107, 8)),6 => std_logic_vector(to_unsigned( 78, 8)),7 => std_logic_vector(to_unsigned( 18, 8)),8 => std_logic_vector(to_unsigned( 72, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 270) then
				RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),1 => std_logic_vector(to_unsigned( 38, 8)),2 => std_logic_vector(to_unsigned( 108, 8)),3 => std_logic_vector(to_unsigned( 80, 8)),4 => std_logic_vector(to_unsigned( 24, 8)),5 => std_logic_vector(to_unsigned( 85, 8)),6 => std_logic_vector(to_unsigned( 96, 8)),7 => std_logic_vector(to_unsigned( 1, 8)),8 => std_logic_vector(to_unsigned( 57, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 271) then
				RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),1 => std_logic_vector(to_unsigned( 62, 8)),2 => std_logic_vector(to_unsigned( 86, 8)),3 => std_logic_vector(to_unsigned( 76, 8)),4 => std_logic_vector(to_unsigned( 21, 8)),5 => std_logic_vector(to_unsigned( 113, 8)),6 => std_logic_vector(to_unsigned( 90, 8)),7 => std_logic_vector(to_unsigned( 124, 8)),8 => std_logic_vector(to_unsigned( 109, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 272) then
				RAM <= (0 => std_logic_vector(to_unsigned( 54, 8)),1 => std_logic_vector(to_unsigned( 9, 8)),2 => std_logic_vector(to_unsigned( 35, 8)),3 => std_logic_vector(to_unsigned( 69, 8)),4 => std_logic_vector(to_unsigned( 46, 8)),5 => std_logic_vector(to_unsigned( 102, 8)),6 => std_logic_vector(to_unsigned( 84, 8)),7 => std_logic_vector(to_unsigned( 107, 8)),8 => std_logic_vector(to_unsigned( 104, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 273) then
				RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),1 => std_logic_vector(to_unsigned( 37, 8)),2 => std_logic_vector(to_unsigned( 106, 8)),3 => std_logic_vector(to_unsigned( 58, 8)),4 => std_logic_vector(to_unsigned( 31, 8)),5 => std_logic_vector(to_unsigned( 95, 8)),6 => std_logic_vector(to_unsigned( 7, 8)),7 => std_logic_vector(to_unsigned( 68, 8)),8 => std_logic_vector(to_unsigned( 105, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 274) then
				RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 55, 8)),3 => std_logic_vector(to_unsigned( 106, 8)),4 => std_logic_vector(to_unsigned( 97, 8)),5 => std_logic_vector(to_unsigned( 87, 8)),6 => std_logic_vector(to_unsigned( 50, 8)),7 => std_logic_vector(to_unsigned( 41, 8)),8 => std_logic_vector(to_unsigned( 26, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 275) then
				RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),1 => std_logic_vector(to_unsigned( 54, 8)),2 => std_logic_vector(to_unsigned( 31, 8)),3 => std_logic_vector(to_unsigned( 41, 8)),4 => std_logic_vector(to_unsigned( 58, 8)),5 => std_logic_vector(to_unsigned( 100, 8)),6 => std_logic_vector(to_unsigned( 5, 8)),7 => std_logic_vector(to_unsigned( 17, 8)),8 => std_logic_vector(to_unsigned( 4, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 276) then
				RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),1 => std_logic_vector(to_unsigned( 84, 8)),2 => std_logic_vector(to_unsigned( 38, 8)),3 => std_logic_vector(to_unsigned( 100, 8)),4 => std_logic_vector(to_unsigned( 105, 8)),5 => std_logic_vector(to_unsigned( 30, 8)),6 => std_logic_vector(to_unsigned( 96, 8)),7 => std_logic_vector(to_unsigned( 13, 8)),8 => std_logic_vector(to_unsigned( 15, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 277) then
				RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),1 => std_logic_vector(to_unsigned( 86, 8)),2 => std_logic_vector(to_unsigned( 51, 8)),3 => std_logic_vector(to_unsigned( 62, 8)),4 => std_logic_vector(to_unsigned( 120, 8)),5 => std_logic_vector(to_unsigned( 73, 8)),6 => std_logic_vector(to_unsigned( 24, 8)),7 => std_logic_vector(to_unsigned( 47, 8)),8 => std_logic_vector(to_unsigned( 125, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 278) then
				RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),1 => std_logic_vector(to_unsigned( 98, 8)),2 => std_logic_vector(to_unsigned( 104, 8)),3 => std_logic_vector(to_unsigned( 51, 8)),4 => std_logic_vector(to_unsigned( 31, 8)),5 => std_logic_vector(to_unsigned( 87, 8)),6 => std_logic_vector(to_unsigned( 94, 8)),7 => std_logic_vector(to_unsigned( 38, 8)),8 => std_logic_vector(to_unsigned( 118, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 279) then
				RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),1 => std_logic_vector(to_unsigned( 83, 8)),2 => std_logic_vector(to_unsigned( 14, 8)),3 => std_logic_vector(to_unsigned( 47, 8)),4 => std_logic_vector(to_unsigned( 94, 8)),5 => std_logic_vector(to_unsigned( 105, 8)),6 => std_logic_vector(to_unsigned( 43, 8)),7 => std_logic_vector(to_unsigned( 31, 8)),8 => std_logic_vector(to_unsigned( 111, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 280) then
				RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),1 => std_logic_vector(to_unsigned( 35, 8)),2 => std_logic_vector(to_unsigned( 16, 8)),3 => std_logic_vector(to_unsigned( 84, 8)),4 => std_logic_vector(to_unsigned( 41, 8)),5 => std_logic_vector(to_unsigned( 62, 8)),6 => std_logic_vector(to_unsigned( 103, 8)),7 => std_logic_vector(to_unsigned( 2, 8)),8 => std_logic_vector(to_unsigned( 74, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 281) then
				RAM <= (0 => std_logic_vector(to_unsigned( 84, 8)),1 => std_logic_vector(to_unsigned( 116, 8)),2 => std_logic_vector(to_unsigned( 72, 8)),3 => std_logic_vector(to_unsigned( 58, 8)),4 => std_logic_vector(to_unsigned( 9, 8)),5 => std_logic_vector(to_unsigned( 35, 8)),6 => std_logic_vector(to_unsigned( 91, 8)),7 => std_logic_vector(to_unsigned( 54, 8)),8 => std_logic_vector(to_unsigned( 118, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 282) then
				RAM <= (0 => std_logic_vector(to_unsigned( 34, 8)),1 => std_logic_vector(to_unsigned( 68, 8)),2 => std_logic_vector(to_unsigned( 88, 8)),3 => std_logic_vector(to_unsigned( 100, 8)),4 => std_logic_vector(to_unsigned( 75, 8)),5 => std_logic_vector(to_unsigned( 40, 8)),6 => std_logic_vector(to_unsigned( 11, 8)),7 => std_logic_vector(to_unsigned( 3, 8)),8 => std_logic_vector(to_unsigned( 47, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 283) then
				RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),1 => std_logic_vector(to_unsigned( 13, 8)),2 => std_logic_vector(to_unsigned( 32, 8)),3 => std_logic_vector(to_unsigned( 97, 8)),4 => std_logic_vector(to_unsigned( 17, 8)),5 => std_logic_vector(to_unsigned( 1, 8)),6 => std_logic_vector(to_unsigned( 65, 8)),7 => std_logic_vector(to_unsigned( 108, 8)),8 => std_logic_vector(to_unsigned( 59, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 284) then
				RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),1 => std_logic_vector(to_unsigned( 112, 8)),2 => std_logic_vector(to_unsigned( 55, 8)),3 => std_logic_vector(to_unsigned( 29, 8)),4 => std_logic_vector(to_unsigned( 119, 8)),5 => std_logic_vector(to_unsigned( 99, 8)),6 => std_logic_vector(to_unsigned( 43, 8)),7 => std_logic_vector(to_unsigned( 20, 8)),8 => std_logic_vector(to_unsigned( 115, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 285) then
				RAM <= (0 => std_logic_vector(to_unsigned( 91, 8)),1 => std_logic_vector(to_unsigned( 36, 8)),2 => std_logic_vector(to_unsigned( 78, 8)),3 => std_logic_vector(to_unsigned( 104, 8)),4 => std_logic_vector(to_unsigned( 18, 8)),5 => std_logic_vector(to_unsigned( 122, 8)),6 => std_logic_vector(to_unsigned( 2, 8)),7 => std_logic_vector(to_unsigned( 8, 8)),8 => std_logic_vector(to_unsigned( 83, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 286) then
				RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),1 => std_logic_vector(to_unsigned( 113, 8)),2 => std_logic_vector(to_unsigned( 59, 8)),3 => std_logic_vector(to_unsigned( 49, 8)),4 => std_logic_vector(to_unsigned( 45, 8)),5 => std_logic_vector(to_unsigned( 63, 8)),6 => std_logic_vector(to_unsigned( 30, 8)),7 => std_logic_vector(to_unsigned( 123, 8)),8 => std_logic_vector(to_unsigned( 116, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 287) then
				RAM <= (0 => std_logic_vector(to_unsigned( 36, 8)),1 => std_logic_vector(to_unsigned( 1, 8)),2 => std_logic_vector(to_unsigned( 52, 8)),3 => std_logic_vector(to_unsigned( 122, 8)),4 => std_logic_vector(to_unsigned( 68, 8)),5 => std_logic_vector(to_unsigned( 7, 8)),6 => std_logic_vector(to_unsigned( 101, 8)),7 => std_logic_vector(to_unsigned( 89, 8)),8 => std_logic_vector(to_unsigned( 42, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 288) then
				RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),1 => std_logic_vector(to_unsigned( 37, 8)),2 => std_logic_vector(to_unsigned( 60, 8)),3 => std_logic_vector(to_unsigned( 86, 8)),4 => std_logic_vector(to_unsigned( 75, 8)),5 => std_logic_vector(to_unsigned( 70, 8)),6 => std_logic_vector(to_unsigned( 64, 8)),7 => std_logic_vector(to_unsigned( 6, 8)),8 => std_logic_vector(to_unsigned( 41, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 289) then
				RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),1 => std_logic_vector(to_unsigned( 81, 8)),2 => std_logic_vector(to_unsigned( 6, 8)),3 => std_logic_vector(to_unsigned( 43, 8)),4 => std_logic_vector(to_unsigned( 91, 8)),5 => std_logic_vector(to_unsigned( 21, 8)),6 => std_logic_vector(to_unsigned( 56, 8)),7 => std_logic_vector(to_unsigned( 38, 8)),8 => std_logic_vector(to_unsigned( 44, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 290) then
				RAM <= (0 => std_logic_vector(to_unsigned( 99, 8)),1 => std_logic_vector(to_unsigned( 112, 8)),2 => std_logic_vector(to_unsigned( 59, 8)),3 => std_logic_vector(to_unsigned( 45, 8)),4 => std_logic_vector(to_unsigned( 52, 8)),5 => std_logic_vector(to_unsigned( 3, 8)),6 => std_logic_vector(to_unsigned( 104, 8)),7 => std_logic_vector(to_unsigned( 69, 8)),8 => std_logic_vector(to_unsigned( 67, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 291) then
				RAM <= (0 => std_logic_vector(to_unsigned( 40, 8)),1 => std_logic_vector(to_unsigned( 28, 8)),2 => std_logic_vector(to_unsigned( 35, 8)),3 => std_logic_vector(to_unsigned( 92, 8)),4 => std_logic_vector(to_unsigned( 83, 8)),5 => std_logic_vector(to_unsigned( 71, 8)),6 => std_logic_vector(to_unsigned( 22, 8)),7 => std_logic_vector(to_unsigned( 116, 8)),8 => std_logic_vector(to_unsigned( 108, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 292) then
				RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),1 => std_logic_vector(to_unsigned( 11, 8)),2 => std_logic_vector(to_unsigned( 116, 8)),3 => std_logic_vector(to_unsigned( 121, 8)),4 => std_logic_vector(to_unsigned( 16, 8)),5 => std_logic_vector(to_unsigned( 102, 8)),6 => std_logic_vector(to_unsigned( 42, 8)),7 => std_logic_vector(to_unsigned( 67, 8)),8 => std_logic_vector(to_unsigned( 43, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 293) then
				RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 85, 8)),3 => std_logic_vector(to_unsigned( 105, 8)),4 => std_logic_vector(to_unsigned( 61, 8)),5 => std_logic_vector(to_unsigned( 2, 8)),6 => std_logic_vector(to_unsigned( 8, 8)),7 => std_logic_vector(to_unsigned( 122, 8)),8 => std_logic_vector(to_unsigned( 34, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 294) then
				RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),1 => std_logic_vector(to_unsigned( 83, 8)),2 => std_logic_vector(to_unsigned( 101, 8)),3 => std_logic_vector(to_unsigned( 109, 8)),4 => std_logic_vector(to_unsigned( 64, 8)),5 => std_logic_vector(to_unsigned( 53, 8)),6 => std_logic_vector(to_unsigned( 32, 8)),7 => std_logic_vector(to_unsigned( 40, 8)),8 => std_logic_vector(to_unsigned( 92, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 295) then
				RAM <= (0 => std_logic_vector(to_unsigned( 110, 8)),1 => std_logic_vector(to_unsigned( 38, 8)),2 => std_logic_vector(to_unsigned( 70, 8)),3 => std_logic_vector(to_unsigned( 47, 8)),4 => std_logic_vector(to_unsigned( 82, 8)),5 => std_logic_vector(to_unsigned( 105, 8)),6 => std_logic_vector(to_unsigned( 11, 8)),7 => std_logic_vector(to_unsigned( 120, 8)),8 => std_logic_vector(to_unsigned( 75, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 296) then
				RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),1 => std_logic_vector(to_unsigned( 81, 8)),2 => std_logic_vector(to_unsigned( 10, 8)),3 => std_logic_vector(to_unsigned( 93, 8)),4 => std_logic_vector(to_unsigned( 118, 8)),5 => std_logic_vector(to_unsigned( 47, 8)),6 => std_logic_vector(to_unsigned( 100, 8)),7 => std_logic_vector(to_unsigned( 54, 8)),8 => std_logic_vector(to_unsigned( 123, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 297) then
				RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),1 => std_logic_vector(to_unsigned( 17, 8)),2 => std_logic_vector(to_unsigned( 5, 8)),3 => std_logic_vector(to_unsigned( 58, 8)),4 => std_logic_vector(to_unsigned( 25, 8)),5 => std_logic_vector(to_unsigned( 97, 8)),6 => std_logic_vector(to_unsigned( 63, 8)),7 => std_logic_vector(to_unsigned( 11, 8)),8 => std_logic_vector(to_unsigned( 83, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 298) then
				RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),1 => std_logic_vector(to_unsigned( 113, 8)),2 => std_logic_vector(to_unsigned( 123, 8)),3 => std_logic_vector(to_unsigned( 4, 8)),4 => std_logic_vector(to_unsigned( 105, 8)),5 => std_logic_vector(to_unsigned( 80, 8)),6 => std_logic_vector(to_unsigned( 76, 8)),7 => std_logic_vector(to_unsigned( 117, 8)),8 => std_logic_vector(to_unsigned( 94, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 299) then
				RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),1 => std_logic_vector(to_unsigned( 123, 8)),2 => std_logic_vector(to_unsigned( 93, 8)),3 => std_logic_vector(to_unsigned( 100, 8)),4 => std_logic_vector(to_unsigned( 20, 8)),5 => std_logic_vector(to_unsigned( 37, 8)),6 => std_logic_vector(to_unsigned( 116, 8)),7 => std_logic_vector(to_unsigned( 26, 8)),8 => std_logic_vector(to_unsigned( 40, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 300) then
				RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),1 => std_logic_vector(to_unsigned( 58, 8)),2 => std_logic_vector(to_unsigned( 32, 8)),3 => std_logic_vector(to_unsigned( 90, 8)),4 => std_logic_vector(to_unsigned( 41, 8)),5 => std_logic_vector(to_unsigned( 115, 8)),6 => std_logic_vector(to_unsigned( 83, 8)),7 => std_logic_vector(to_unsigned( 76, 8)),8 => std_logic_vector(to_unsigned( 56, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 301) then
				RAM <= (0 => std_logic_vector(to_unsigned( 107, 8)),1 => std_logic_vector(to_unsigned( 6, 8)),2 => std_logic_vector(to_unsigned( 39, 8)),3 => std_logic_vector(to_unsigned( 50, 8)),4 => std_logic_vector(to_unsigned( 0, 8)),5 => std_logic_vector(to_unsigned( 15, 8)),6 => std_logic_vector(to_unsigned( 99, 8)),7 => std_logic_vector(to_unsigned( 94, 8)),8 => std_logic_vector(to_unsigned( 1, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 302) then
				RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),1 => std_logic_vector(to_unsigned( 123, 8)),2 => std_logic_vector(to_unsigned( 100, 8)),3 => std_logic_vector(to_unsigned( 54, 8)),4 => std_logic_vector(to_unsigned( 47, 8)),5 => std_logic_vector(to_unsigned( 116, 8)),6 => std_logic_vector(to_unsigned( 0, 8)),7 => std_logic_vector(to_unsigned( 31, 8)),8 => std_logic_vector(to_unsigned( 111, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 303) then
				RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 54, 8)),3 => std_logic_vector(to_unsigned( 82, 8)),4 => std_logic_vector(to_unsigned( 77, 8)),5 => std_logic_vector(to_unsigned( 107, 8)),6 => std_logic_vector(to_unsigned( 33, 8)),7 => std_logic_vector(to_unsigned( 92, 8)),8 => std_logic_vector(to_unsigned( 59, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 304) then
				RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),1 => std_logic_vector(to_unsigned( 28, 8)),2 => std_logic_vector(to_unsigned( 70, 8)),3 => std_logic_vector(to_unsigned( 51, 8)),4 => std_logic_vector(to_unsigned( 44, 8)),5 => std_logic_vector(to_unsigned( 109, 8)),6 => std_logic_vector(to_unsigned( 6, 8)),7 => std_logic_vector(to_unsigned( 90, 8)),8 => std_logic_vector(to_unsigned( 68, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 305) then
				RAM <= (0 => std_logic_vector(to_unsigned( 25, 8)),1 => std_logic_vector(to_unsigned( 17, 8)),2 => std_logic_vector(to_unsigned( 1, 8)),3 => std_logic_vector(to_unsigned( 79, 8)),4 => std_logic_vector(to_unsigned( 83, 8)),5 => std_logic_vector(to_unsigned( 34, 8)),6 => std_logic_vector(to_unsigned( 73, 8)),7 => std_logic_vector(to_unsigned( 61, 8)),8 => std_logic_vector(to_unsigned( 55, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 306) then
				RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),1 => std_logic_vector(to_unsigned( 119, 8)),2 => std_logic_vector(to_unsigned( 96, 8)),3 => std_logic_vector(to_unsigned( 115, 8)),4 => std_logic_vector(to_unsigned( 102, 8)),5 => std_logic_vector(to_unsigned( 34, 8)),6 => std_logic_vector(to_unsigned( 3, 8)),7 => std_logic_vector(to_unsigned( 49, 8)),8 => std_logic_vector(to_unsigned( 52, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 307) then
				RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),1 => std_logic_vector(to_unsigned( 19, 8)),2 => std_logic_vector(to_unsigned( 71, 8)),3 => std_logic_vector(to_unsigned( 4, 8)),4 => std_logic_vector(to_unsigned( 32, 8)),5 => std_logic_vector(to_unsigned( 41, 8)),6 => std_logic_vector(to_unsigned( 110, 8)),7 => std_logic_vector(to_unsigned( 8, 8)),8 => std_logic_vector(to_unsigned( 54, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 308) then
				RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),1 => std_logic_vector(to_unsigned( 102, 8)),2 => std_logic_vector(to_unsigned( 15, 8)),3 => std_logic_vector(to_unsigned( 74, 8)),4 => std_logic_vector(to_unsigned( 6, 8)),5 => std_logic_vector(to_unsigned( 38, 8)),6 => std_logic_vector(to_unsigned( 48, 8)),7 => std_logic_vector(to_unsigned( 95, 8)),8 => std_logic_vector(to_unsigned( 35, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 309) then
				RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),1 => std_logic_vector(to_unsigned( 44, 8)),2 => std_logic_vector(to_unsigned( 100, 8)),3 => std_logic_vector(to_unsigned( 122, 8)),4 => std_logic_vector(to_unsigned( 82, 8)),5 => std_logic_vector(to_unsigned( 58, 8)),6 => std_logic_vector(to_unsigned( 20, 8)),7 => std_logic_vector(to_unsigned( 93, 8)),8 => std_logic_vector(to_unsigned( 63, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 310) then
				RAM <= (0 => std_logic_vector(to_unsigned( 9, 8)),1 => std_logic_vector(to_unsigned( 116, 8)),2 => std_logic_vector(to_unsigned( 34, 8)),3 => std_logic_vector(to_unsigned( 20, 8)),4 => std_logic_vector(to_unsigned( 65, 8)),5 => std_logic_vector(to_unsigned( 53, 8)),6 => std_logic_vector(to_unsigned( 98, 8)),7 => std_logic_vector(to_unsigned( 92, 8)),8 => std_logic_vector(to_unsigned( 120, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 311) then
				RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),1 => std_logic_vector(to_unsigned( 7, 8)),2 => std_logic_vector(to_unsigned( 61, 8)),3 => std_logic_vector(to_unsigned( 87, 8)),4 => std_logic_vector(to_unsigned( 52, 8)),5 => std_logic_vector(to_unsigned( 67, 8)),6 => std_logic_vector(to_unsigned( 113, 8)),7 => std_logic_vector(to_unsigned( 40, 8)),8 => std_logic_vector(to_unsigned( 97, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 312) then
				RAM <= (0 => std_logic_vector(to_unsigned( 61, 8)),1 => std_logic_vector(to_unsigned( 114, 8)),2 => std_logic_vector(to_unsigned( 89, 8)),3 => std_logic_vector(to_unsigned( 32, 8)),4 => std_logic_vector(to_unsigned( 48, 8)),5 => std_logic_vector(to_unsigned( 8, 8)),6 => std_logic_vector(to_unsigned( 99, 8)),7 => std_logic_vector(to_unsigned( 105, 8)),8 => std_logic_vector(to_unsigned( 90, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 313) then
				RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),1 => std_logic_vector(to_unsigned( 119, 8)),2 => std_logic_vector(to_unsigned( 63, 8)),3 => std_logic_vector(to_unsigned( 115, 8)),4 => std_logic_vector(to_unsigned( 23, 8)),5 => std_logic_vector(to_unsigned( 101, 8)),6 => std_logic_vector(to_unsigned( 91, 8)),7 => std_logic_vector(to_unsigned( 80, 8)),8 => std_logic_vector(to_unsigned( 59, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 314) then
				RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),1 => std_logic_vector(to_unsigned( 94, 8)),2 => std_logic_vector(to_unsigned( 123, 8)),3 => std_logic_vector(to_unsigned( 26, 8)),4 => std_logic_vector(to_unsigned( 64, 8)),5 => std_logic_vector(to_unsigned( 42, 8)),6 => std_logic_vector(to_unsigned( 68, 8)),7 => std_logic_vector(to_unsigned( 30, 8)),8 => std_logic_vector(to_unsigned( 39, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 315) then
				RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),1 => std_logic_vector(to_unsigned( 57, 8)),2 => std_logic_vector(to_unsigned( 99, 8)),3 => std_logic_vector(to_unsigned( 119, 8)),4 => std_logic_vector(to_unsigned( 44, 8)),5 => std_logic_vector(to_unsigned( 64, 8)),6 => std_logic_vector(to_unsigned( 33, 8)),7 => std_logic_vector(to_unsigned( 6, 8)),8 => std_logic_vector(to_unsigned( 29, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 316) then
				RAM <= (0 => std_logic_vector(to_unsigned( 112, 8)),1 => std_logic_vector(to_unsigned( 20, 8)),2 => std_logic_vector(to_unsigned( 45, 8)),3 => std_logic_vector(to_unsigned( 14, 8)),4 => std_logic_vector(to_unsigned( 60, 8)),5 => std_logic_vector(to_unsigned( 32, 8)),6 => std_logic_vector(to_unsigned( 25, 8)),7 => std_logic_vector(to_unsigned( 55, 8)),8 => std_logic_vector(to_unsigned( 92, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 317) then
				RAM <= (0 => std_logic_vector(to_unsigned( 11, 8)),1 => std_logic_vector(to_unsigned( 102, 8)),2 => std_logic_vector(to_unsigned( 22, 8)),3 => std_logic_vector(to_unsigned( 95, 8)),4 => std_logic_vector(to_unsigned( 113, 8)),5 => std_logic_vector(to_unsigned( 87, 8)),6 => std_logic_vector(to_unsigned( 38, 8)),7 => std_logic_vector(to_unsigned( 75, 8)),8 => std_logic_vector(to_unsigned( 61, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 318) then
				RAM <= (0 => std_logic_vector(to_unsigned( 84, 8)),1 => std_logic_vector(to_unsigned( 40, 8)),2 => std_logic_vector(to_unsigned( 123, 8)),3 => std_logic_vector(to_unsigned( 47, 8)),4 => std_logic_vector(to_unsigned( 88, 8)),5 => std_logic_vector(to_unsigned( 14, 8)),6 => std_logic_vector(to_unsigned( 0, 8)),7 => std_logic_vector(to_unsigned( 6, 8)),8 => std_logic_vector(to_unsigned( 21, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 319) then
				RAM <= (0 => std_logic_vector(to_unsigned( 12, 8)),1 => std_logic_vector(to_unsigned( 54, 8)),2 => std_logic_vector(to_unsigned( 63, 8)),3 => std_logic_vector(to_unsigned( 107, 8)),4 => std_logic_vector(to_unsigned( 34, 8)),5 => std_logic_vector(to_unsigned( 42, 8)),6 => std_logic_vector(to_unsigned( 97, 8)),7 => std_logic_vector(to_unsigned( 80, 8)),8 => std_logic_vector(to_unsigned( 109, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 320) then
				RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),1 => std_logic_vector(to_unsigned( 36, 8)),2 => std_logic_vector(to_unsigned( 16, 8)),3 => std_logic_vector(to_unsigned( 32, 8)),4 => std_logic_vector(to_unsigned( 84, 8)),5 => std_logic_vector(to_unsigned( 59, 8)),6 => std_logic_vector(to_unsigned( 100, 8)),7 => std_logic_vector(to_unsigned( 76, 8)),8 => std_logic_vector(to_unsigned( 111, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 321) then
				RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),1 => std_logic_vector(to_unsigned( 6, 8)),2 => std_logic_vector(to_unsigned( 26, 8)),3 => std_logic_vector(to_unsigned( 81, 8)),4 => std_logic_vector(to_unsigned( 1, 8)),5 => std_logic_vector(to_unsigned( 17, 8)),6 => std_logic_vector(to_unsigned( 89, 8)),7 => std_logic_vector(to_unsigned( 44, 8)),8 => std_logic_vector(to_unsigned( 62, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 322) then
				RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),1 => std_logic_vector(to_unsigned( 5, 8)),2 => std_logic_vector(to_unsigned( 29, 8)),3 => std_logic_vector(to_unsigned( 25, 8)),4 => std_logic_vector(to_unsigned( 96, 8)),5 => std_logic_vector(to_unsigned( 83, 8)),6 => std_logic_vector(to_unsigned( 55, 8)),7 => std_logic_vector(to_unsigned( 78, 8)),8 => std_logic_vector(to_unsigned( 8, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 323) then
				RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),1 => std_logic_vector(to_unsigned( 100, 8)),2 => std_logic_vector(to_unsigned( 67, 8)),3 => std_logic_vector(to_unsigned( 2, 8)),4 => std_logic_vector(to_unsigned( 58, 8)),5 => std_logic_vector(to_unsigned( 26, 8)),6 => std_logic_vector(to_unsigned( 116, 8)),7 => std_logic_vector(to_unsigned( 42, 8)),8 => std_logic_vector(to_unsigned( 38, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 324) then
				RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),1 => std_logic_vector(to_unsigned( 25, 8)),2 => std_logic_vector(to_unsigned( 0, 8)),3 => std_logic_vector(to_unsigned( 113, 8)),4 => std_logic_vector(to_unsigned( 36, 8)),5 => std_logic_vector(to_unsigned( 107, 8)),6 => std_logic_vector(to_unsigned( 58, 8)),7 => std_logic_vector(to_unsigned( 90, 8)),8 => std_logic_vector(to_unsigned( 72, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 325) then
				RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),1 => std_logic_vector(to_unsigned( 40, 8)),2 => std_logic_vector(to_unsigned( 33, 8)),3 => std_logic_vector(to_unsigned( 89, 8)),4 => std_logic_vector(to_unsigned( 117, 8)),5 => std_logic_vector(to_unsigned( 82, 8)),6 => std_logic_vector(to_unsigned( 20, 8)),7 => std_logic_vector(to_unsigned( 103, 8)),8 => std_logic_vector(to_unsigned( 49, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 326) then
				RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),1 => std_logic_vector(to_unsigned( 78, 8)),2 => std_logic_vector(to_unsigned( 91, 8)),3 => std_logic_vector(to_unsigned( 15, 8)),4 => std_logic_vector(to_unsigned( 107, 8)),5 => std_logic_vector(to_unsigned( 70, 8)),6 => std_logic_vector(to_unsigned( 9, 8)),7 => std_logic_vector(to_unsigned( 39, 8)),8 => std_logic_vector(to_unsigned( 36, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 327) then
				RAM <= (0 => std_logic_vector(to_unsigned( 119, 8)),1 => std_logic_vector(to_unsigned( 109, 8)),2 => std_logic_vector(to_unsigned( 19, 8)),3 => std_logic_vector(to_unsigned( 94, 8)),4 => std_logic_vector(to_unsigned( 80, 8)),5 => std_logic_vector(to_unsigned( 64, 8)),6 => std_logic_vector(to_unsigned( 115, 8)),7 => std_logic_vector(to_unsigned( 51, 8)),8 => std_logic_vector(to_unsigned( 79, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 328) then
				RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),1 => std_logic_vector(to_unsigned( 123, 8)),2 => std_logic_vector(to_unsigned( 33, 8)),3 => std_logic_vector(to_unsigned( 29, 8)),4 => std_logic_vector(to_unsigned( 115, 8)),5 => std_logic_vector(to_unsigned( 47, 8)),6 => std_logic_vector(to_unsigned( 109, 8)),7 => std_logic_vector(to_unsigned( 101, 8)),8 => std_logic_vector(to_unsigned( 92, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 329) then
				RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),1 => std_logic_vector(to_unsigned( 51, 8)),2 => std_logic_vector(to_unsigned( 116, 8)),3 => std_logic_vector(to_unsigned( 100, 8)),4 => std_logic_vector(to_unsigned( 91, 8)),5 => std_logic_vector(to_unsigned( 105, 8)),6 => std_logic_vector(to_unsigned( 21, 8)),7 => std_logic_vector(to_unsigned( 74, 8)),8 => std_logic_vector(to_unsigned( 112, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 330) then
				RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),1 => std_logic_vector(to_unsigned( 48, 8)),2 => std_logic_vector(to_unsigned( 117, 8)),3 => std_logic_vector(to_unsigned( 89, 8)),4 => std_logic_vector(to_unsigned( 2, 8)),5 => std_logic_vector(to_unsigned( 41, 8)),6 => std_logic_vector(to_unsigned( 13, 8)),7 => std_logic_vector(to_unsigned( 7, 8)),8 => std_logic_vector(to_unsigned( 111, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 331) then
				RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),1 => std_logic_vector(to_unsigned( 65, 8)),2 => std_logic_vector(to_unsigned( 15, 8)),3 => std_logic_vector(to_unsigned( 11, 8)),4 => std_logic_vector(to_unsigned( 94, 8)),5 => std_logic_vector(to_unsigned( 26, 8)),6 => std_logic_vector(to_unsigned( 56, 8)),7 => std_logic_vector(to_unsigned( 111, 8)),8 => std_logic_vector(to_unsigned( 65, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 332) then
				RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 25, 8)),3 => std_logic_vector(to_unsigned( 21, 8)),4 => std_logic_vector(to_unsigned( 80, 8)),5 => std_logic_vector(to_unsigned( 41, 8)),6 => std_logic_vector(to_unsigned( 12, 8)),7 => std_logic_vector(to_unsigned( 88, 8)),8 => std_logic_vector(to_unsigned( 49, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 333) then
				RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),1 => std_logic_vector(to_unsigned( 99, 8)),2 => std_logic_vector(to_unsigned( 91, 8)),3 => std_logic_vector(to_unsigned( 106, 8)),4 => std_logic_vector(to_unsigned( 11, 8)),5 => std_logic_vector(to_unsigned( 51, 8)),6 => std_logic_vector(to_unsigned( 77, 8)),7 => std_logic_vector(to_unsigned( 60, 8)),8 => std_logic_vector(to_unsigned( 126, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 334) then
				RAM <= (0 => std_logic_vector(to_unsigned( 117, 8)),1 => std_logic_vector(to_unsigned( 15, 8)),2 => std_logic_vector(to_unsigned( 106, 8)),3 => std_logic_vector(to_unsigned( 75, 8)),4 => std_logic_vector(to_unsigned( 61, 8)),5 => std_logic_vector(to_unsigned( 97, 8)),6 => std_logic_vector(to_unsigned( 23, 8)),7 => std_logic_vector(to_unsigned( 44, 8)),8 => std_logic_vector(to_unsigned( 59, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 335) then
				RAM <= (0 => std_logic_vector(to_unsigned( 115, 8)),1 => std_logic_vector(to_unsigned( 4, 8)),2 => std_logic_vector(to_unsigned( 47, 8)),3 => std_logic_vector(to_unsigned( 69, 8)),4 => std_logic_vector(to_unsigned( 8, 8)),5 => std_logic_vector(to_unsigned( 97, 8)),6 => std_logic_vector(to_unsigned( 80, 8)),7 => std_logic_vector(to_unsigned( 64, 8)),8 => std_logic_vector(to_unsigned( 87, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 336) then
				RAM <= (0 => std_logic_vector(to_unsigned( 60, 8)),1 => std_logic_vector(to_unsigned( 118, 8)),2 => std_logic_vector(to_unsigned( 45, 8)),3 => std_logic_vector(to_unsigned( 11, 8)),4 => std_logic_vector(to_unsigned( 109, 8)),5 => std_logic_vector(to_unsigned( 64, 8)),6 => std_logic_vector(to_unsigned( 93, 8)),7 => std_logic_vector(to_unsigned( 75, 8)),8 => std_logic_vector(to_unsigned( 100, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 337) then
				RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),1 => std_logic_vector(to_unsigned( 84, 8)),2 => std_logic_vector(to_unsigned( 107, 8)),3 => std_logic_vector(to_unsigned( 100, 8)),4 => std_logic_vector(to_unsigned( 64, 8)),5 => std_logic_vector(to_unsigned( 27, 8)),6 => std_logic_vector(to_unsigned( 4, 8)),7 => std_logic_vector(to_unsigned( 59, 8)),8 => std_logic_vector(to_unsigned( 50, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 338) then
				RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),1 => std_logic_vector(to_unsigned( 77, 8)),2 => std_logic_vector(to_unsigned( 67, 8)),3 => std_logic_vector(to_unsigned( 9, 8)),4 => std_logic_vector(to_unsigned( 95, 8)),5 => std_logic_vector(to_unsigned( 54, 8)),6 => std_logic_vector(to_unsigned( 48, 8)),7 => std_logic_vector(to_unsigned( 42, 8)),8 => std_logic_vector(to_unsigned( 79, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 339) then
				RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),1 => std_logic_vector(to_unsigned( 7, 8)),2 => std_logic_vector(to_unsigned( 49, 8)),3 => std_logic_vector(to_unsigned( 19, 8)),4 => std_logic_vector(to_unsigned( 106, 8)),5 => std_logic_vector(to_unsigned( 86, 8)),6 => std_logic_vector(to_unsigned( 59, 8)),7 => std_logic_vector(to_unsigned( 102, 8)),8 => std_logic_vector(to_unsigned( 29, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 340) then
				RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),1 => std_logic_vector(to_unsigned( 26, 8)),2 => std_logic_vector(to_unsigned( 123, 8)),3 => std_logic_vector(to_unsigned( 119, 8)),4 => std_logic_vector(to_unsigned( 2, 8)),5 => std_logic_vector(to_unsigned( 47, 8)),6 => std_logic_vector(to_unsigned( 60, 8)),7 => std_logic_vector(to_unsigned( 41, 8)),8 => std_logic_vector(to_unsigned( 71, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 341) then
				RAM <= (0 => std_logic_vector(to_unsigned( 45, 8)),1 => std_logic_vector(to_unsigned( 100, 8)),2 => std_logic_vector(to_unsigned( 34, 8)),3 => std_logic_vector(to_unsigned( 119, 8)),4 => std_logic_vector(to_unsigned( 73, 8)),5 => std_logic_vector(to_unsigned( 5, 8)),6 => std_logic_vector(to_unsigned( 12, 8)),7 => std_logic_vector(to_unsigned( 112, 8)),8 => std_logic_vector(to_unsigned( 124, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 342) then
				RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),1 => std_logic_vector(to_unsigned( 13, 8)),2 => std_logic_vector(to_unsigned( 32, 8)),3 => std_logic_vector(to_unsigned( 107, 8)),4 => std_logic_vector(to_unsigned( 73, 8)),5 => std_logic_vector(to_unsigned( 91, 8)),6 => std_logic_vector(to_unsigned( 54, 8)),7 => std_logic_vector(to_unsigned( 101, 8)),8 => std_logic_vector(to_unsigned( 89, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 343) then
				RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),1 => std_logic_vector(to_unsigned( 32, 8)),2 => std_logic_vector(to_unsigned( 55, 8)),3 => std_logic_vector(to_unsigned( 74, 8)),4 => std_logic_vector(to_unsigned( 110, 8)),5 => std_logic_vector(to_unsigned( 114, 8)),6 => std_logic_vector(to_unsigned( 100, 8)),7 => std_logic_vector(to_unsigned( 80, 8)),8 => std_logic_vector(to_unsigned( 77, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 344) then
				RAM <= (0 => std_logic_vector(to_unsigned( 103, 8)),1 => std_logic_vector(to_unsigned( 7, 8)),2 => std_logic_vector(to_unsigned( 29, 8)),3 => std_logic_vector(to_unsigned( 65, 8)),4 => std_logic_vector(to_unsigned( 12, 8)),5 => std_logic_vector(to_unsigned( 97, 8)),6 => std_logic_vector(to_unsigned( 61, 8)),7 => std_logic_vector(to_unsigned( 3, 8)),8 => std_logic_vector(to_unsigned( 22, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 345) then
				RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),1 => std_logic_vector(to_unsigned( 37, 8)),2 => std_logic_vector(to_unsigned( 112, 8)),3 => std_logic_vector(to_unsigned( 83, 8)),4 => std_logic_vector(to_unsigned( 117, 8)),5 => std_logic_vector(to_unsigned( 67, 8)),6 => std_logic_vector(to_unsigned( 88, 8)),7 => std_logic_vector(to_unsigned( 59, 8)),8 => std_logic_vector(to_unsigned( 21, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 346) then
				RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),1 => std_logic_vector(to_unsigned( 65, 8)),2 => std_logic_vector(to_unsigned( 82, 8)),3 => std_logic_vector(to_unsigned( 120, 8)),4 => std_logic_vector(to_unsigned( 115, 8)),5 => std_logic_vector(to_unsigned( 31, 8)),6 => std_logic_vector(to_unsigned( 12, 8)),7 => std_logic_vector(to_unsigned( 96, 8)),8 => std_logic_vector(to_unsigned( 82, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 347) then
				RAM <= (0 => std_logic_vector(to_unsigned( 100, 8)),1 => std_logic_vector(to_unsigned( 20, 8)),2 => std_logic_vector(to_unsigned( 90, 8)),3 => std_logic_vector(to_unsigned( 76, 8)),4 => std_logic_vector(to_unsigned( 42, 8)),5 => std_logic_vector(to_unsigned( 6, 8)),6 => std_logic_vector(to_unsigned( 25, 8)),7 => std_logic_vector(to_unsigned( 71, 8)),8 => std_logic_vector(to_unsigned( 78, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 348) then
				RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),1 => std_logic_vector(to_unsigned( 1, 8)),2 => std_logic_vector(to_unsigned( 8, 8)),3 => std_logic_vector(to_unsigned( 30, 8)),4 => std_logic_vector(to_unsigned( 112, 8)),5 => std_logic_vector(to_unsigned( 75, 8)),6 => std_logic_vector(to_unsigned( 16, 8)),7 => std_logic_vector(to_unsigned( 38, 8)),8 => std_logic_vector(to_unsigned( 28, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 349) then
				RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),1 => std_logic_vector(to_unsigned( 115, 8)),2 => std_logic_vector(to_unsigned( 64, 8)),3 => std_logic_vector(to_unsigned( 2, 8)),4 => std_logic_vector(to_unsigned( 29, 8)),5 => std_logic_vector(to_unsigned( 91, 8)),6 => std_logic_vector(to_unsigned( 25, 8)),7 => std_logic_vector(to_unsigned( 83, 8)),8 => std_logic_vector(to_unsigned( 34, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 350) then
				RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),1 => std_logic_vector(to_unsigned( 92, 8)),2 => std_logic_vector(to_unsigned( 105, 8)),3 => std_logic_vector(to_unsigned( 30, 8)),4 => std_logic_vector(to_unsigned( 63, 8)),5 => std_logic_vector(to_unsigned( 69, 8)),6 => std_logic_vector(to_unsigned( 35, 8)),7 => std_logic_vector(to_unsigned( 111, 8)),8 => std_logic_vector(to_unsigned( 124, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 351) then
				RAM <= (0 => std_logic_vector(to_unsigned( 20, 8)),1 => std_logic_vector(to_unsigned( 107, 8)),2 => std_logic_vector(to_unsigned( 82, 8)),3 => std_logic_vector(to_unsigned( 99, 8)),4 => std_logic_vector(to_unsigned( 9, 8)),5 => std_logic_vector(to_unsigned( 38, 8)),6 => std_logic_vector(to_unsigned( 50, 8)),7 => std_logic_vector(to_unsigned( 64, 8)),8 => std_logic_vector(to_unsigned( 33, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 352) then
				RAM <= (0 => std_logic_vector(to_unsigned( 65, 8)),1 => std_logic_vector(to_unsigned( 14, 8)),2 => std_logic_vector(to_unsigned( 36, 8)),3 => std_logic_vector(to_unsigned( 31, 8)),4 => std_logic_vector(to_unsigned( 46, 8)),5 => std_logic_vector(to_unsigned( 110, 8)),6 => std_logic_vector(to_unsigned( 73, 8)),7 => std_logic_vector(to_unsigned( 4, 8)),8 => std_logic_vector(to_unsigned( 9, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 353) then
				RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),1 => std_logic_vector(to_unsigned( 120, 8)),2 => std_logic_vector(to_unsigned( 59, 8)),3 => std_logic_vector(to_unsigned( 69, 8)),4 => std_logic_vector(to_unsigned( 47, 8)),5 => std_logic_vector(to_unsigned( 16, 8)),6 => std_logic_vector(to_unsigned( 83, 8)),7 => std_logic_vector(to_unsigned( 7, 8)),8 => std_logic_vector(to_unsigned( 59, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 354) then
				RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),1 => std_logic_vector(to_unsigned( 1, 8)),2 => std_logic_vector(to_unsigned( 47, 8)),3 => std_logic_vector(to_unsigned( 85, 8)),4 => std_logic_vector(to_unsigned( 123, 8)),5 => std_logic_vector(to_unsigned( 74, 8)),6 => std_logic_vector(to_unsigned( 14, 8)),7 => std_logic_vector(to_unsigned( 20, 8)),8 => std_logic_vector(to_unsigned( 72, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 355) then
				RAM <= (0 => std_logic_vector(to_unsigned( 22, 8)),1 => std_logic_vector(to_unsigned( 93, 8)),2 => std_logic_vector(to_unsigned( 59, 8)),3 => std_logic_vector(to_unsigned( 50, 8)),4 => std_logic_vector(to_unsigned( 65, 8)),5 => std_logic_vector(to_unsigned( 73, 8)),6 => std_logic_vector(to_unsigned( 86, 8)),7 => std_logic_vector(to_unsigned( 15, 8)),8 => std_logic_vector(to_unsigned( 72, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 356) then
				RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),1 => std_logic_vector(to_unsigned( 46, 8)),2 => std_logic_vector(to_unsigned( 124, 8)),3 => std_logic_vector(to_unsigned( 63, 8)),4 => std_logic_vector(to_unsigned( 110, 8)),5 => std_logic_vector(to_unsigned( 119, 8)),6 => std_logic_vector(to_unsigned( 35, 8)),7 => std_logic_vector(to_unsigned( 101, 8)),8 => std_logic_vector(to_unsigned( 9, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 357) then
				RAM <= (0 => std_logic_vector(to_unsigned( 13, 8)),1 => std_logic_vector(to_unsigned( 76, 8)),2 => std_logic_vector(to_unsigned( 121, 8)),3 => std_logic_vector(to_unsigned( 47, 8)),4 => std_logic_vector(to_unsigned( 4, 8)),5 => std_logic_vector(to_unsigned( 26, 8)),6 => std_logic_vector(to_unsigned( 112, 8)),7 => std_logic_vector(to_unsigned( 92, 8)),8 => std_logic_vector(to_unsigned( 79, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 358) then
				RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),1 => std_logic_vector(to_unsigned( 45, 8)),2 => std_logic_vector(to_unsigned( 107, 8)),3 => std_logic_vector(to_unsigned( 16, 8)),4 => std_logic_vector(to_unsigned( 20, 8)),5 => std_logic_vector(to_unsigned( 101, 8)),6 => std_logic_vector(to_unsigned( 85, 8)),7 => std_logic_vector(to_unsigned( 26, 8)),8 => std_logic_vector(to_unsigned( 73, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 359) then
				RAM <= (0 => std_logic_vector(to_unsigned( 91, 8)),1 => std_logic_vector(to_unsigned( 63, 8)),2 => std_logic_vector(to_unsigned( 48, 8)),3 => std_logic_vector(to_unsigned( 52, 8)),4 => std_logic_vector(to_unsigned( 1, 8)),5 => std_logic_vector(to_unsigned( 30, 8)),6 => std_logic_vector(to_unsigned( 107, 8)),7 => std_logic_vector(to_unsigned( 7, 8)),8 => std_logic_vector(to_unsigned( 31, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 360) then
				RAM <= (0 => std_logic_vector(to_unsigned( 106, 8)),1 => std_logic_vector(to_unsigned( 82, 8)),2 => std_logic_vector(to_unsigned( 50, 8)),3 => std_logic_vector(to_unsigned( 89, 8)),4 => std_logic_vector(to_unsigned( 101, 8)),5 => std_logic_vector(to_unsigned( 58, 8)),6 => std_logic_vector(to_unsigned( 77, 8)),7 => std_logic_vector(to_unsigned( 38, 8)),8 => std_logic_vector(to_unsigned( 5, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 361) then
				RAM <= (0 => std_logic_vector(to_unsigned( 46, 8)),1 => std_logic_vector(to_unsigned( 50, 8)),2 => std_logic_vector(to_unsigned( 55, 8)),3 => std_logic_vector(to_unsigned( 12, 8)),4 => std_logic_vector(to_unsigned( 7, 8)),5 => std_logic_vector(to_unsigned( 25, 8)),6 => std_logic_vector(to_unsigned( 112, 8)),7 => std_logic_vector(to_unsigned( 34, 8)),8 => std_logic_vector(to_unsigned( 31, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 362) then
				RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),1 => std_logic_vector(to_unsigned( 23, 8)),2 => std_logic_vector(to_unsigned( 109, 8)),3 => std_logic_vector(to_unsigned( 45, 8)),4 => std_logic_vector(to_unsigned( 76, 8)),5 => std_logic_vector(to_unsigned( 39, 8)),6 => std_logic_vector(to_unsigned( 65, 8)),7 => std_logic_vector(to_unsigned( 14, 8)),8 => std_logic_vector(to_unsigned( 116, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 363) then
				RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),1 => std_logic_vector(to_unsigned( 124, 8)),2 => std_logic_vector(to_unsigned( 35, 8)),3 => std_logic_vector(to_unsigned( 58, 8)),4 => std_logic_vector(to_unsigned( 65, 8)),5 => std_logic_vector(to_unsigned( 18, 8)),6 => std_logic_vector(to_unsigned( 111, 8)),7 => std_logic_vector(to_unsigned( 80, 8)),8 => std_logic_vector(to_unsigned( 110, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 364) then
				RAM <= (0 => std_logic_vector(to_unsigned( 94, 8)),1 => std_logic_vector(to_unsigned( 81, 8)),2 => std_logic_vector(to_unsigned( 72, 8)),3 => std_logic_vector(to_unsigned( 113, 8)),4 => std_logic_vector(to_unsigned( 118, 8)),5 => std_logic_vector(to_unsigned( 23, 8)),6 => std_logic_vector(to_unsigned( 76, 8)),7 => std_logic_vector(to_unsigned( 18, 8)),8 => std_logic_vector(to_unsigned( 27, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 365) then
				RAM <= (0 => std_logic_vector(to_unsigned( 42, 8)),1 => std_logic_vector(to_unsigned( 85, 8)),2 => std_logic_vector(to_unsigned( 103, 8)),3 => std_logic_vector(to_unsigned( 37, 8)),4 => std_logic_vector(to_unsigned( 117, 8)),5 => std_logic_vector(to_unsigned( 65, 8)),6 => std_logic_vector(to_unsigned( 89, 8)),7 => std_logic_vector(to_unsigned( 58, 8)),8 => std_logic_vector(to_unsigned( 125, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 366) then
				RAM <= (0 => std_logic_vector(to_unsigned( 30, 8)),1 => std_logic_vector(to_unsigned( 51, 8)),2 => std_logic_vector(to_unsigned( 36, 8)),3 => std_logic_vector(to_unsigned( 95, 8)),4 => std_logic_vector(to_unsigned( 24, 8)),5 => std_logic_vector(to_unsigned( 63, 8)),6 => std_logic_vector(to_unsigned( 87, 8)),7 => std_logic_vector(to_unsigned( 6, 8)),8 => std_logic_vector(to_unsigned( 32, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 367) then
				RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),1 => std_logic_vector(to_unsigned( 68, 8)),2 => std_logic_vector(to_unsigned( 108, 8)),3 => std_logic_vector(to_unsigned( 35, 8)),4 => std_logic_vector(to_unsigned( 121, 8)),5 => std_logic_vector(to_unsigned( 16, 8)),6 => std_logic_vector(to_unsigned( 115, 8)),7 => std_logic_vector(to_unsigned( 90, 8)),8 => std_logic_vector(to_unsigned( 90, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 368) then
				RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),1 => std_logic_vector(to_unsigned( 95, 8)),2 => std_logic_vector(to_unsigned( 62, 8)),3 => std_logic_vector(to_unsigned( 105, 8)),4 => std_logic_vector(to_unsigned( 48, 8)),5 => std_logic_vector(to_unsigned( 9, 8)),6 => std_logic_vector(to_unsigned( 57, 8)),7 => std_logic_vector(to_unsigned( 15, 8)),8 => std_logic_vector(to_unsigned( 95, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 369) then
				RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),1 => std_logic_vector(to_unsigned( 105, 8)),2 => std_logic_vector(to_unsigned( 35, 8)),3 => std_logic_vector(to_unsigned( 59, 8)),4 => std_logic_vector(to_unsigned( 23, 8)),5 => std_logic_vector(to_unsigned( 45, 8)),6 => std_logic_vector(to_unsigned( 93, 8)),7 => std_logic_vector(to_unsigned( 66, 8)),8 => std_logic_vector(to_unsigned( 83, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 370) then
				RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),1 => std_logic_vector(to_unsigned( 44, 8)),2 => std_logic_vector(to_unsigned( 99, 8)),3 => std_logic_vector(to_unsigned( 15, 8)),4 => std_logic_vector(to_unsigned( 2, 8)),5 => std_logic_vector(to_unsigned( 60, 8)),6 => std_logic_vector(to_unsigned( 117, 8)),7 => std_logic_vector(to_unsigned( 95, 8)),8 => std_logic_vector(to_unsigned( 10, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 371) then
				RAM <= (0 => std_logic_vector(to_unsigned( 89, 8)),1 => std_logic_vector(to_unsigned( 4, 8)),2 => std_logic_vector(to_unsigned( 32, 8)),3 => std_logic_vector(to_unsigned( 22, 8)),4 => std_logic_vector(to_unsigned( 83, 8)),5 => std_logic_vector(to_unsigned( 101, 8)),6 => std_logic_vector(to_unsigned( 114, 8)),7 => std_logic_vector(to_unsigned( 44, 8)),8 => std_logic_vector(to_unsigned( 31, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 372) then
				RAM <= (0 => std_logic_vector(to_unsigned( 112, 8)),1 => std_logic_vector(to_unsigned( 65, 8)),2 => std_logic_vector(to_unsigned( 9, 8)),3 => std_logic_vector(to_unsigned( 32, 8)),4 => std_logic_vector(to_unsigned( 58, 8)),5 => std_logic_vector(to_unsigned( 40, 8)),6 => std_logic_vector(to_unsigned( 27, 8)),7 => std_logic_vector(to_unsigned( 18, 8)),8 => std_logic_vector(to_unsigned( 11, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 373) then
				RAM <= (0 => std_logic_vector(to_unsigned( 98, 8)),1 => std_logic_vector(to_unsigned( 85, 8)),2 => std_logic_vector(to_unsigned( 26, 8)),3 => std_logic_vector(to_unsigned( 102, 8)),4 => std_logic_vector(to_unsigned( 45, 8)),5 => std_logic_vector(to_unsigned( 94, 8)),6 => std_logic_vector(to_unsigned( 14, 8)),7 => std_logic_vector(to_unsigned( 119, 8)),8 => std_logic_vector(to_unsigned( 82, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 374) then
				RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),1 => std_logic_vector(to_unsigned( 7, 8)),2 => std_logic_vector(to_unsigned( 99, 8)),3 => std_logic_vector(to_unsigned( 75, 8)),4 => std_logic_vector(to_unsigned( 22, 8)),5 => std_logic_vector(to_unsigned( 104, 8)),6 => std_logic_vector(to_unsigned( 118, 8)),7 => std_logic_vector(to_unsigned( 18, 8)),8 => std_logic_vector(to_unsigned( 61, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 375) then
				RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),1 => std_logic_vector(to_unsigned( 57, 8)),2 => std_logic_vector(to_unsigned( 23, 8)),3 => std_logic_vector(to_unsigned( 85, 8)),4 => std_logic_vector(to_unsigned( 43, 8)),5 => std_logic_vector(to_unsigned( 73, 8)),6 => std_logic_vector(to_unsigned( 18, 8)),7 => std_logic_vector(to_unsigned( 94, 8)),8 => std_logic_vector(to_unsigned( 36, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 376) then
				RAM <= (0 => std_logic_vector(to_unsigned( 55, 8)),1 => std_logic_vector(to_unsigned( 63, 8)),2 => std_logic_vector(to_unsigned( 29, 8)),3 => std_logic_vector(to_unsigned( 106, 8)),4 => std_logic_vector(to_unsigned( 11, 8)),5 => std_logic_vector(to_unsigned( 85, 8)),6 => std_logic_vector(to_unsigned( 90, 8)),7 => std_logic_vector(to_unsigned( 15, 8)),8 => std_logic_vector(to_unsigned( 8, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 377) then
				RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),1 => std_logic_vector(to_unsigned( 70, 8)),2 => std_logic_vector(to_unsigned( 113, 8)),3 => std_logic_vector(to_unsigned( 34, 8)),4 => std_logic_vector(to_unsigned( 24, 8)),5 => std_logic_vector(to_unsigned( 87, 8)),6 => std_logic_vector(to_unsigned( 98, 8)),7 => std_logic_vector(to_unsigned( 104, 8)),8 => std_logic_vector(to_unsigned( 113, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 378) then
				RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),1 => std_logic_vector(to_unsigned( 120, 8)),2 => std_logic_vector(to_unsigned( 11, 8)),3 => std_logic_vector(to_unsigned( 74, 8)),4 => std_logic_vector(to_unsigned( 20, 8)),5 => std_logic_vector(to_unsigned( 2, 8)),6 => std_logic_vector(to_unsigned( 41, 8)),7 => std_logic_vector(to_unsigned( 91, 8)),8 => std_logic_vector(to_unsigned( 110, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 379) then
				RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),1 => std_logic_vector(to_unsigned( 109, 8)),2 => std_logic_vector(to_unsigned( 3, 8)),3 => std_logic_vector(to_unsigned( 71, 8)),4 => std_logic_vector(to_unsigned( 88, 8)),5 => std_logic_vector(to_unsigned( 122, 8)),6 => std_logic_vector(to_unsigned( 16, 8)),7 => std_logic_vector(to_unsigned( 100, 8)),8 => std_logic_vector(to_unsigned( 108, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 380) then
				RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),1 => std_logic_vector(to_unsigned( 52, 8)),2 => std_logic_vector(to_unsigned( 116, 8)),3 => std_logic_vector(to_unsigned( 120, 8)),4 => std_logic_vector(to_unsigned( 93, 8)),5 => std_logic_vector(to_unsigned( 43, 8)),6 => std_logic_vector(to_unsigned( 124, 8)),7 => std_logic_vector(to_unsigned( 12, 8)),8 => std_logic_vector(to_unsigned( 29, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 381) then
				RAM <= (0 => std_logic_vector(to_unsigned( 35, 8)),1 => std_logic_vector(to_unsigned( 29, 8)),2 => std_logic_vector(to_unsigned( 48, 8)),3 => std_logic_vector(to_unsigned( 87, 8)),4 => std_logic_vector(to_unsigned( 72, 8)),5 => std_logic_vector(to_unsigned( 18, 8)),6 => std_logic_vector(to_unsigned( 94, 8)),7 => std_logic_vector(to_unsigned( 77, 8)),8 => std_logic_vector(to_unsigned( 113, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 382) then
				RAM <= (0 => std_logic_vector(to_unsigned( 46, 8)),1 => std_logic_vector(to_unsigned( 19, 8)),2 => std_logic_vector(to_unsigned( 113, 8)),3 => std_logic_vector(to_unsigned( 123, 8)),4 => std_logic_vector(to_unsigned( 117, 8)),5 => std_logic_vector(to_unsigned( 86, 8)),6 => std_logic_vector(to_unsigned( 13, 8)),7 => std_logic_vector(to_unsigned( 97, 8)),8 => std_logic_vector(to_unsigned( 19, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 383) then
				RAM <= (0 => std_logic_vector(to_unsigned( 123, 8)),1 => std_logic_vector(to_unsigned( 59, 8)),2 => std_logic_vector(to_unsigned( 73, 8)),3 => std_logic_vector(to_unsigned( 42, 8)),4 => std_logic_vector(to_unsigned( 77, 8)),5 => std_logic_vector(to_unsigned( 95, 8)),6 => std_logic_vector(to_unsigned( 13, 8)),7 => std_logic_vector(to_unsigned( 21, 8)),8 => std_logic_vector(to_unsigned( 42, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 384) then
				RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),1 => std_logic_vector(to_unsigned( 3, 8)),2 => std_logic_vector(to_unsigned( 105, 8)),3 => std_logic_vector(to_unsigned( 84, 8)),4 => std_logic_vector(to_unsigned( 92, 8)),5 => std_logic_vector(to_unsigned( 64, 8)),6 => std_logic_vector(to_unsigned( 98, 8)),7 => std_logic_vector(to_unsigned( 115, 8)),8 => std_logic_vector(to_unsigned( 4, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 385) then
				RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),1 => std_logic_vector(to_unsigned( 7, 8)),2 => std_logic_vector(to_unsigned( 37, 8)),3 => std_logic_vector(to_unsigned( 90, 8)),4 => std_logic_vector(to_unsigned( 60, 8)),5 => std_logic_vector(to_unsigned( 72, 8)),6 => std_logic_vector(to_unsigned( 2, 8)),7 => std_logic_vector(to_unsigned( 98, 8)),8 => std_logic_vector(to_unsigned( 35, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 386) then
				RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),1 => std_logic_vector(to_unsigned( 102, 8)),2 => std_logic_vector(to_unsigned( 36, 8)),3 => std_logic_vector(to_unsigned( 5, 8)),4 => std_logic_vector(to_unsigned( 118, 8)),5 => std_logic_vector(to_unsigned( 108, 8)),6 => std_logic_vector(to_unsigned( 49, 8)),7 => std_logic_vector(to_unsigned( 30, 8)),8 => std_logic_vector(to_unsigned( 26, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 387) then
				RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),1 => std_logic_vector(to_unsigned( 13, 8)),2 => std_logic_vector(to_unsigned( 111, 8)),3 => std_logic_vector(to_unsigned( 53, 8)),4 => std_logic_vector(to_unsigned( 61, 8)),5 => std_logic_vector(to_unsigned( 32, 8)),6 => std_logic_vector(to_unsigned( 4, 8)),7 => std_logic_vector(to_unsigned( 100, 8)),8 => std_logic_vector(to_unsigned( 46, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 388) then
				RAM <= (0 => std_logic_vector(to_unsigned( 33, 8)),1 => std_logic_vector(to_unsigned( 79, 8)),2 => std_logic_vector(to_unsigned( 105, 8)),3 => std_logic_vector(to_unsigned( 12, 8)),4 => std_logic_vector(to_unsigned( 3, 8)),5 => std_logic_vector(to_unsigned( 115, 8)),6 => std_logic_vector(to_unsigned( 89, 8)),7 => std_logic_vector(to_unsigned( 71, 8)),8 => std_logic_vector(to_unsigned( 127, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 389) then
				RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),1 => std_logic_vector(to_unsigned( 54, 8)),2 => std_logic_vector(to_unsigned( 96, 8)),3 => std_logic_vector(to_unsigned( 91, 8)),4 => std_logic_vector(to_unsigned( 36, 8)),5 => std_logic_vector(to_unsigned( 20, 8)),6 => std_logic_vector(to_unsigned( 48, 8)),7 => std_logic_vector(to_unsigned( 7, 8)),8 => std_logic_vector(to_unsigned( 95, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 390) then
				RAM <= (0 => std_logic_vector(to_unsigned( 51, 8)),1 => std_logic_vector(to_unsigned( 5, 8)),2 => std_logic_vector(to_unsigned( 116, 8)),3 => std_logic_vector(to_unsigned( 41, 8)),4 => std_logic_vector(to_unsigned( 76, 8)),5 => std_logic_vector(to_unsigned( 1, 8)),6 => std_logic_vector(to_unsigned( 55, 8)),7 => std_logic_vector(to_unsigned( 98, 8)),8 => std_logic_vector(to_unsigned( 116, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 391) then
				RAM <= (0 => std_logic_vector(to_unsigned( 8, 8)),1 => std_logic_vector(to_unsigned( 120, 8)),2 => std_logic_vector(to_unsigned( 124, 8)),3 => std_logic_vector(to_unsigned( 57, 8)),4 => std_logic_vector(to_unsigned( 21, 8)),5 => std_logic_vector(to_unsigned( 31, 8)),6 => std_logic_vector(to_unsigned( 106, 8)),7 => std_logic_vector(to_unsigned( 97, 8)),8 => std_logic_vector(to_unsigned( 40, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 392) then
				RAM <= (0 => std_logic_vector(to_unsigned( 88, 8)),1 => std_logic_vector(to_unsigned( 7, 8)),2 => std_logic_vector(to_unsigned( 94, 8)),3 => std_logic_vector(to_unsigned( 112, 8)),4 => std_logic_vector(to_unsigned( 81, 8)),5 => std_logic_vector(to_unsigned( 43, 8)),6 => std_logic_vector(to_unsigned( 2, 8)),7 => std_logic_vector(to_unsigned( 62, 8)),8 => std_logic_vector(to_unsigned( 86, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 393) then
				RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),1 => std_logic_vector(to_unsigned( 31, 8)),2 => std_logic_vector(to_unsigned( 78, 8)),3 => std_logic_vector(to_unsigned( 66, 8)),4 => std_logic_vector(to_unsigned( 107, 8)),5 => std_logic_vector(to_unsigned( 57, 8)),6 => std_logic_vector(to_unsigned( 51, 8)),7 => std_logic_vector(to_unsigned( 114, 8)),8 => std_logic_vector(to_unsigned( 13, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 394) then
				RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),1 => std_logic_vector(to_unsigned( 110, 8)),2 => std_logic_vector(to_unsigned( 94, 8)),3 => std_logic_vector(to_unsigned( 99, 8)),4 => std_logic_vector(to_unsigned( 51, 8)),5 => std_logic_vector(to_unsigned( 45, 8)),6 => std_logic_vector(to_unsigned( 24, 8)),7 => std_logic_vector(to_unsigned( 6, 8)),8 => std_logic_vector(to_unsigned( 24, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 395) then
				RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),1 => std_logic_vector(to_unsigned( 98, 8)),2 => std_logic_vector(to_unsigned( 108, 8)),3 => std_logic_vector(to_unsigned( 90, 8)),4 => std_logic_vector(to_unsigned( 35, 8)),5 => std_logic_vector(to_unsigned( 16, 8)),6 => std_logic_vector(to_unsigned( 44, 8)),7 => std_logic_vector(to_unsigned( 29, 8)),8 => std_logic_vector(to_unsigned( 8, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 396) then
				RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),1 => std_logic_vector(to_unsigned( 49, 8)),2 => std_logic_vector(to_unsigned( 121, 8)),3 => std_logic_vector(to_unsigned( 64, 8)),4 => std_logic_vector(to_unsigned( 80, 8)),5 => std_logic_vector(to_unsigned( 117, 8)),6 => std_logic_vector(to_unsigned( 97, 8)),7 => std_logic_vector(to_unsigned( 88, 8)),8 => std_logic_vector(to_unsigned( 25, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 397) then
				RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),1 => std_logic_vector(to_unsigned( 40, 8)),2 => std_logic_vector(to_unsigned( 83, 8)),3 => std_logic_vector(to_unsigned( 90, 8)),4 => std_logic_vector(to_unsigned( 19, 8)),5 => std_logic_vector(to_unsigned( 107, 8)),6 => std_logic_vector(to_unsigned( 98, 8)),7 => std_logic_vector(to_unsigned( 30, 8)),8 => std_logic_vector(to_unsigned( 120, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 398) then
				RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),1 => std_logic_vector(to_unsigned( 65, 8)),2 => std_logic_vector(to_unsigned( 89, 8)),3 => std_logic_vector(to_unsigned( 19, 8)),4 => std_logic_vector(to_unsigned( 31, 8)),5 => std_logic_vector(to_unsigned( 110, 8)),6 => std_logic_vector(to_unsigned( 78, 8)),7 => std_logic_vector(to_unsigned( 3, 8)),8 => std_logic_vector(to_unsigned( 5, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 399) then
				RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),1 => std_logic_vector(to_unsigned( 29, 8)),2 => std_logic_vector(to_unsigned( 41, 8)),3 => std_logic_vector(to_unsigned( 46, 8)),4 => std_logic_vector(to_unsigned( 86, 8)),5 => std_logic_vector(to_unsigned( 68, 8)),6 => std_logic_vector(to_unsigned( 59, 8)),7 => std_logic_vector(to_unsigned( 64, 8)),8 => std_logic_vector(to_unsigned( 90, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 400) then
				RAM <= (0 => std_logic_vector(to_unsigned( 72, 8)),1 => std_logic_vector(to_unsigned( 123, 8)),2 => std_logic_vector(to_unsigned( 11, 8)),3 => std_logic_vector(to_unsigned( 82, 8)),4 => std_logic_vector(to_unsigned( 55, 8)),5 => std_logic_vector(to_unsigned( 33, 8)),6 => std_logic_vector(to_unsigned( 67, 8)),7 => std_logic_vector(to_unsigned( 42, 8)),8 => std_logic_vector(to_unsigned( 29, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 401) then
				RAM <= (0 => std_logic_vector(to_unsigned( 8, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 31, 8)),3 => std_logic_vector(to_unsigned( 13, 8)),4 => std_logic_vector(to_unsigned( 18, 8)),5 => std_logic_vector(to_unsigned( 41, 8)),6 => std_logic_vector(to_unsigned( 49, 8)),7 => std_logic_vector(to_unsigned( 111, 8)),8 => std_logic_vector(to_unsigned( 50, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 402) then
				RAM <= (0 => std_logic_vector(to_unsigned( 74, 8)),1 => std_logic_vector(to_unsigned( 57, 8)),2 => std_logic_vector(to_unsigned( 100, 8)),3 => std_logic_vector(to_unsigned( 49, 8)),4 => std_logic_vector(to_unsigned( 85, 8)),5 => std_logic_vector(to_unsigned( 3, 8)),6 => std_logic_vector(to_unsigned( 7, 8)),7 => std_logic_vector(to_unsigned( 114, 8)),8 => std_logic_vector(to_unsigned( 75, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 403) then
				RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),1 => std_logic_vector(to_unsigned( 1, 8)),2 => std_logic_vector(to_unsigned( 41, 8)),3 => std_logic_vector(to_unsigned( 85, 8)),4 => std_logic_vector(to_unsigned( 55, 8)),5 => std_logic_vector(to_unsigned( 103, 8)),6 => std_logic_vector(to_unsigned( 121, 8)),7 => std_logic_vector(to_unsigned( 61, 8)),8 => std_logic_vector(to_unsigned( 103, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 404) then
				RAM <= (0 => std_logic_vector(to_unsigned( 68, 8)),1 => std_logic_vector(to_unsigned( 49, 8)),2 => std_logic_vector(to_unsigned( 73, 8)),3 => std_logic_vector(to_unsigned( 121, 8)),4 => std_logic_vector(to_unsigned( 90, 8)),5 => std_logic_vector(to_unsigned( 25, 8)),6 => std_logic_vector(to_unsigned( 94, 8)),7 => std_logic_vector(to_unsigned( 83, 8)),8 => std_logic_vector(to_unsigned( 107, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 405) then
				RAM <= (0 => std_logic_vector(to_unsigned( 57, 8)),1 => std_logic_vector(to_unsigned( 12, 8)),2 => std_logic_vector(to_unsigned( 83, 8)),3 => std_logic_vector(to_unsigned( 109, 8)),4 => std_logic_vector(to_unsigned( 68, 8)),5 => std_logic_vector(to_unsigned( 17, 8)),6 => std_logic_vector(to_unsigned( 89, 8)),7 => std_logic_vector(to_unsigned( 47, 8)),8 => std_logic_vector(to_unsigned( 32, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 406) then
				RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),1 => std_logic_vector(to_unsigned( 93, 8)),2 => std_logic_vector(to_unsigned( 86, 8)),3 => std_logic_vector(to_unsigned( 109, 8)),4 => std_logic_vector(to_unsigned( 115, 8)),5 => std_logic_vector(to_unsigned( 47, 8)),6 => std_logic_vector(to_unsigned( 26, 8)),7 => std_logic_vector(to_unsigned( 3, 8)),8 => std_logic_vector(to_unsigned( 85, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 407) then
				RAM <= (0 => std_logic_vector(to_unsigned( 79, 8)),1 => std_logic_vector(to_unsigned( 15, 8)),2 => std_logic_vector(to_unsigned( 29, 8)),3 => std_logic_vector(to_unsigned( 108, 8)),4 => std_logic_vector(to_unsigned( 57, 8)),5 => std_logic_vector(to_unsigned( 1, 8)),6 => std_logic_vector(to_unsigned( 39, 8)),7 => std_logic_vector(to_unsigned( 48, 8)),8 => std_logic_vector(to_unsigned( 118, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 408) then
				RAM <= (0 => std_logic_vector(to_unsigned( 49, 8)),1 => std_logic_vector(to_unsigned( 20, 8)),2 => std_logic_vector(to_unsigned( 42, 8)),3 => std_logic_vector(to_unsigned( 29, 8)),4 => std_logic_vector(to_unsigned( 12, 8)),5 => std_logic_vector(to_unsigned( 93, 8)),6 => std_logic_vector(to_unsigned( 38, 8)),7 => std_logic_vector(to_unsigned( 110, 8)),8 => std_logic_vector(to_unsigned( 45, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 409) then
				RAM <= (0 => std_logic_vector(to_unsigned( 43, 8)),1 => std_logic_vector(to_unsigned( 122, 8)),2 => std_logic_vector(to_unsigned( 71, 8)),3 => std_logic_vector(to_unsigned( 7, 8)),4 => std_logic_vector(to_unsigned( 48, 8)),5 => std_logic_vector(to_unsigned( 21, 8)),6 => std_logic_vector(to_unsigned( 56, 8)),7 => std_logic_vector(to_unsigned( 92, 8)),8 => std_logic_vector(to_unsigned( 43, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 410) then
				RAM <= (0 => std_logic_vector(to_unsigned( 42, 8)),1 => std_logic_vector(to_unsigned( 25, 8)),2 => std_logic_vector(to_unsigned( 103, 8)),3 => std_logic_vector(to_unsigned( 53, 8)),4 => std_logic_vector(to_unsigned( 77, 8)),5 => std_logic_vector(to_unsigned( 72, 8)),6 => std_logic_vector(to_unsigned( 93, 8)),7 => std_logic_vector(to_unsigned( 121, 8)),8 => std_logic_vector(to_unsigned( 54, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 411) then
				RAM <= (0 => std_logic_vector(to_unsigned( 76, 8)),1 => std_logic_vector(to_unsigned( 101, 8)),2 => std_logic_vector(to_unsigned( 27, 8)),3 => std_logic_vector(to_unsigned( 4, 8)),4 => std_logic_vector(to_unsigned( 116, 8)),5 => std_logic_vector(to_unsigned( 72, 8)),6 => std_logic_vector(to_unsigned( 66, 8)),7 => std_logic_vector(to_unsigned( 97, 8)),8 => std_logic_vector(to_unsigned( 61, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 412) then
				RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),1 => std_logic_vector(to_unsigned( 42, 8)),2 => std_logic_vector(to_unsigned( 37, 8)),3 => std_logic_vector(to_unsigned( 115, 8)),4 => std_logic_vector(to_unsigned( 7, 8)),5 => std_logic_vector(to_unsigned( 19, 8)),6 => std_logic_vector(to_unsigned( 104, 8)),7 => std_logic_vector(to_unsigned( 32, 8)),8 => std_logic_vector(to_unsigned( 85, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 413) then
				RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),1 => std_logic_vector(to_unsigned( 120, 8)),2 => std_logic_vector(to_unsigned( 102, 8)),3 => std_logic_vector(to_unsigned( 8, 8)),4 => std_logic_vector(to_unsigned( 31, 8)),5 => std_logic_vector(to_unsigned( 54, 8)),6 => std_logic_vector(to_unsigned( 37, 8)),7 => std_logic_vector(to_unsigned( 69, 8)),8 => std_logic_vector(to_unsigned( 78, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 414) then
				RAM <= (0 => std_logic_vector(to_unsigned( 53, 8)),1 => std_logic_vector(to_unsigned( 109, 8)),2 => std_logic_vector(to_unsigned( 48, 8)),3 => std_logic_vector(to_unsigned( 90, 8)),4 => std_logic_vector(to_unsigned( 17, 8)),5 => std_logic_vector(to_unsigned( 84, 8)),6 => std_logic_vector(to_unsigned( 11, 8)),7 => std_logic_vector(to_unsigned( 0, 8)),8 => std_logic_vector(to_unsigned( 60, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 415) then
				RAM <= (0 => std_logic_vector(to_unsigned( 78, 8)),1 => std_logic_vector(to_unsigned( 47, 8)),2 => std_logic_vector(to_unsigned( 37, 8)),3 => std_logic_vector(to_unsigned( 29, 8)),4 => std_logic_vector(to_unsigned( 83, 8)),5 => std_logic_vector(to_unsigned( 114, 8)),6 => std_logic_vector(to_unsigned( 120, 8)),7 => std_logic_vector(to_unsigned( 7, 8)),8 => std_logic_vector(to_unsigned( 4, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 416) then
				RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),1 => std_logic_vector(to_unsigned( 92, 8)),2 => std_logic_vector(to_unsigned( 106, 8)),3 => std_logic_vector(to_unsigned( 79, 8)),4 => std_logic_vector(to_unsigned( 50, 8)),5 => std_logic_vector(to_unsigned( 15, 8)),6 => std_logic_vector(to_unsigned( 7, 8)),7 => std_logic_vector(to_unsigned( 117, 8)),8 => std_logic_vector(to_unsigned( 26, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 417) then
				RAM <= (0 => std_logic_vector(to_unsigned( 16, 8)),1 => std_logic_vector(to_unsigned( 96, 8)),2 => std_logic_vector(to_unsigned( 28, 8)),3 => std_logic_vector(to_unsigned( 11, 8)),4 => std_logic_vector(to_unsigned( 36, 8)),5 => std_logic_vector(to_unsigned( 69, 8)),6 => std_logic_vector(to_unsigned( 49, 8)),7 => std_logic_vector(to_unsigned( 61, 8)),8 => std_logic_vector(to_unsigned( 121, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 418) then
				RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),1 => std_logic_vector(to_unsigned( 76, 8)),2 => std_logic_vector(to_unsigned( 21, 8)),3 => std_logic_vector(to_unsigned( 100, 8)),4 => std_logic_vector(to_unsigned( 10, 8)),5 => std_logic_vector(to_unsigned( 94, 8)),6 => std_logic_vector(to_unsigned( 25, 8)),7 => std_logic_vector(to_unsigned( 81, 8)),8 => std_logic_vector(to_unsigned( 57, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 419) then
				RAM <= (0 => std_logic_vector(to_unsigned( 46, 8)),1 => std_logic_vector(to_unsigned( 101, 8)),2 => std_logic_vector(to_unsigned( 79, 8)),3 => std_logic_vector(to_unsigned( 117, 8)),4 => std_logic_vector(to_unsigned( 107, 8)),5 => std_logic_vector(to_unsigned( 56, 8)),6 => std_logic_vector(to_unsigned( 84, 8)),7 => std_logic_vector(to_unsigned( 35, 8)),8 => std_logic_vector(to_unsigned( 17, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 420) then
				RAM <= (0 => std_logic_vector(to_unsigned( 104, 8)),1 => std_logic_vector(to_unsigned( 50, 8)),2 => std_logic_vector(to_unsigned( 35, 8)),3 => std_logic_vector(to_unsigned( 108, 8)),4 => std_logic_vector(to_unsigned( 10, 8)),5 => std_logic_vector(to_unsigned( 6, 8)),6 => std_logic_vector(to_unsigned( 87, 8)),7 => std_logic_vector(to_unsigned( 124, 8)),8 => std_logic_vector(to_unsigned( 27, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 421) then
				RAM <= (0 => std_logic_vector(to_unsigned( 19, 8)),1 => std_logic_vector(to_unsigned( 31, 8)),2 => std_logic_vector(to_unsigned( 75, 8)),3 => std_logic_vector(to_unsigned( 14, 8)),4 => std_logic_vector(to_unsigned( 100, 8)),5 => std_logic_vector(to_unsigned( 82, 8)),6 => std_logic_vector(to_unsigned( 44, 8)),7 => std_logic_vector(to_unsigned( 94, 8)),8 => std_logic_vector(to_unsigned( 0, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 422) then
				RAM <= (0 => std_logic_vector(to_unsigned( 97, 8)),1 => std_logic_vector(to_unsigned( 60, 8)),2 => std_logic_vector(to_unsigned( 115, 8)),3 => std_logic_vector(to_unsigned( 5, 8)),4 => std_logic_vector(to_unsigned( 103, 8)),5 => std_logic_vector(to_unsigned( 14, 8)),6 => std_logic_vector(to_unsigned( 28, 8)),7 => std_logic_vector(to_unsigned( 78, 8)),8 => std_logic_vector(to_unsigned( 51, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 423) then
				RAM <= (0 => std_logic_vector(to_unsigned( 21, 8)),1 => std_logic_vector(to_unsigned( 14, 8)),2 => std_logic_vector(to_unsigned( 0, 8)),3 => std_logic_vector(to_unsigned( 40, 8)),4 => std_logic_vector(to_unsigned( 30, 8)),5 => std_logic_vector(to_unsigned( 59, 8)),6 => std_logic_vector(to_unsigned( 93, 8)),7 => std_logic_vector(to_unsigned( 85, 8)),8 => std_logic_vector(to_unsigned( 117, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 424) then
				RAM <= (0 => std_logic_vector(to_unsigned( 95, 8)),1 => std_logic_vector(to_unsigned( 27, 8)),2 => std_logic_vector(to_unsigned( 112, 8)),3 => std_logic_vector(to_unsigned( 62, 8)),4 => std_logic_vector(to_unsigned( 2, 8)),5 => std_logic_vector(to_unsigned( 15, 8)),6 => std_logic_vector(to_unsigned( 70, 8)),7 => std_logic_vector(to_unsigned( 31, 8)),8 => std_logic_vector(to_unsigned( 16, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 425) then
				RAM <= (0 => std_logic_vector(to_unsigned( 91, 8)),1 => std_logic_vector(to_unsigned( 52, 8)),2 => std_logic_vector(to_unsigned( 102, 8)),3 => std_logic_vector(to_unsigned( 21, 8)),4 => std_logic_vector(to_unsigned( 124, 8)),5 => std_logic_vector(to_unsigned( 35, 8)),6 => std_logic_vector(to_unsigned( 109, 8)),7 => std_logic_vector(to_unsigned( 86, 8)),8 => std_logic_vector(to_unsigned( 42, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 426) then
				RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),1 => std_logic_vector(to_unsigned( 59, 8)),2 => std_logic_vector(to_unsigned( 25, 8)),3 => std_logic_vector(to_unsigned( 97, 8)),4 => std_logic_vector(to_unsigned( 16, 8)),5 => std_logic_vector(to_unsigned( 87, 8)),6 => std_logic_vector(to_unsigned( 83, 8)),7 => std_logic_vector(to_unsigned( 8, 8)),8 => std_logic_vector(to_unsigned( 96, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 427) then
				RAM <= (0 => std_logic_vector(to_unsigned( 80, 8)),1 => std_logic_vector(to_unsigned( 46, 8)),2 => std_logic_vector(to_unsigned( 14, 8)),3 => std_logic_vector(to_unsigned( 57, 8)),4 => std_logic_vector(to_unsigned( 31, 8)),5 => std_logic_vector(to_unsigned( 95, 8)),6 => std_logic_vector(to_unsigned( 120, 8)),7 => std_logic_vector(to_unsigned( 6, 8)),8 => std_logic_vector(to_unsigned( 76, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 428) then
				RAM <= (0 => std_logic_vector(to_unsigned( 101, 8)),1 => std_logic_vector(to_unsigned( 70, 8)),2 => std_logic_vector(to_unsigned( 81, 8)),3 => std_logic_vector(to_unsigned( 0, 8)),4 => std_logic_vector(to_unsigned( 39, 8)),5 => std_logic_vector(to_unsigned( 52, 8)),6 => std_logic_vector(to_unsigned( 26, 8)),7 => std_logic_vector(to_unsigned( 66, 8)),8 => std_logic_vector(to_unsigned( 46, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 429) then
				RAM <= (0 => std_logic_vector(to_unsigned( 102, 8)),1 => std_logic_vector(to_unsigned( 29, 8)),2 => std_logic_vector(to_unsigned( 47, 8)),3 => std_logic_vector(to_unsigned( 37, 8)),4 => std_logic_vector(to_unsigned( 62, 8)),5 => std_logic_vector(to_unsigned( 119, 8)),6 => std_logic_vector(to_unsigned( 33, 8)),7 => std_logic_vector(to_unsigned( 83, 8)),8 => std_logic_vector(to_unsigned( 117, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 430) then
				RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),1 => std_logic_vector(to_unsigned( 18, 8)),2 => std_logic_vector(to_unsigned( 75, 8)),3 => std_logic_vector(to_unsigned( 10, 8)),4 => std_logic_vector(to_unsigned( 59, 8)),5 => std_logic_vector(to_unsigned( 105, 8)),6 => std_logic_vector(to_unsigned( 111, 8)),7 => std_logic_vector(to_unsigned( 43, 8)),8 => std_logic_vector(to_unsigned( 114, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 431) then
				RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),1 => std_logic_vector(to_unsigned( 72, 8)),2 => std_logic_vector(to_unsigned( 106, 8)),3 => std_logic_vector(to_unsigned( 113, 8)),4 => std_logic_vector(to_unsigned( 12, 8)),5 => std_logic_vector(to_unsigned( 23, 8)),6 => std_logic_vector(to_unsigned( 16, 8)),7 => std_logic_vector(to_unsigned( 50, 8)),8 => std_logic_vector(to_unsigned( 77, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 432) then
				RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),1 => std_logic_vector(to_unsigned( 41, 8)),2 => std_logic_vector(to_unsigned( 7, 8)),3 => std_logic_vector(to_unsigned( 56, 8)),4 => std_logic_vector(to_unsigned( 89, 8)),5 => std_logic_vector(to_unsigned( 30, 8)),6 => std_logic_vector(to_unsigned( 76, 8)),7 => std_logic_vector(to_unsigned( 81, 8)),8 => std_logic_vector(to_unsigned( 12, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 433) then
				RAM <= (0 => std_logic_vector(to_unsigned( 85, 8)),1 => std_logic_vector(to_unsigned( 40, 8)),2 => std_logic_vector(to_unsigned( 77, 8)),3 => std_logic_vector(to_unsigned( 25, 8)),4 => std_logic_vector(to_unsigned( 110, 8)),5 => std_logic_vector(to_unsigned( 51, 8)),6 => std_logic_vector(to_unsigned( 94, 8)),7 => std_logic_vector(to_unsigned( 69, 8)),8 => std_logic_vector(to_unsigned( 76, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 434) then
				RAM <= (0 => std_logic_vector(to_unsigned( 52, 8)),1 => std_logic_vector(to_unsigned( 0, 8)),2 => std_logic_vector(to_unsigned( 8, 8)),3 => std_logic_vector(to_unsigned( 107, 8)),4 => std_logic_vector(to_unsigned( 36, 8)),5 => std_logic_vector(to_unsigned( 82, 8)),6 => std_logic_vector(to_unsigned( 93, 8)),7 => std_logic_vector(to_unsigned( 69, 8)),8 => std_logic_vector(to_unsigned( 117, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 435) then
				RAM <= (0 => std_logic_vector(to_unsigned( 42, 8)),1 => std_logic_vector(to_unsigned( 5, 8)),2 => std_logic_vector(to_unsigned( 76, 8)),3 => std_logic_vector(to_unsigned( 65, 8)),4 => std_logic_vector(to_unsigned( 80, 8)),5 => std_logic_vector(to_unsigned( 57, 8)),6 => std_logic_vector(to_unsigned( 112, 8)),7 => std_logic_vector(to_unsigned( 53, 8)),8 => std_logic_vector(to_unsigned( 77, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 436) then
				RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),1 => std_logic_vector(to_unsigned( 23, 8)),2 => std_logic_vector(to_unsigned( 78, 8)),3 => std_logic_vector(to_unsigned( 61, 8)),4 => std_logic_vector(to_unsigned( 87, 8)),5 => std_logic_vector(to_unsigned( 57, 8)),6 => std_logic_vector(to_unsigned( 47, 8)),7 => std_logic_vector(to_unsigned( 51, 8)),8 => std_logic_vector(to_unsigned( 118, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 437) then
				RAM <= (0 => std_logic_vector(to_unsigned( 7, 8)),1 => std_logic_vector(to_unsigned( 103, 8)),2 => std_logic_vector(to_unsigned( 30, 8)),3 => std_logic_vector(to_unsigned( 72, 8)),4 => std_logic_vector(to_unsigned( 67, 8)),5 => std_logic_vector(to_unsigned( 47, 8)),6 => std_logic_vector(to_unsigned( 12, 8)),7 => std_logic_vector(to_unsigned( 122, 8)),8 => std_logic_vector(to_unsigned( 45, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 438) then
				RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),1 => std_logic_vector(to_unsigned( 101, 8)),2 => std_logic_vector(to_unsigned( 112, 8)),3 => std_logic_vector(to_unsigned( 41, 8)),4 => std_logic_vector(to_unsigned( 88, 8)),5 => std_logic_vector(to_unsigned( 20, 8)),6 => std_logic_vector(to_unsigned( 124, 8)),7 => std_logic_vector(to_unsigned( 59, 8)),8 => std_logic_vector(to_unsigned( 126, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 439) then
				RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),1 => std_logic_vector(to_unsigned( 86, 8)),2 => std_logic_vector(to_unsigned( 115, 8)),3 => std_logic_vector(to_unsigned( 98, 8)),4 => std_logic_vector(to_unsigned( 57, 8)),5 => std_logic_vector(to_unsigned( 66, 8)),6 => std_logic_vector(to_unsigned( 78, 8)),7 => std_logic_vector(to_unsigned( 110, 8)),8 => std_logic_vector(to_unsigned( 56, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 440) then
				RAM <= (0 => std_logic_vector(to_unsigned( 24, 8)),1 => std_logic_vector(to_unsigned( 71, 8)),2 => std_logic_vector(to_unsigned( 118, 8)),3 => std_logic_vector(to_unsigned( 47, 8)),4 => std_logic_vector(to_unsigned( 38, 8)),5 => std_logic_vector(to_unsigned( 8, 8)),6 => std_logic_vector(to_unsigned( 95, 8)),7 => std_logic_vector(to_unsigned( 104, 8)),8 => std_logic_vector(to_unsigned( 125, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 441) then
				RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),1 => std_logic_vector(to_unsigned( 49, 8)),2 => std_logic_vector(to_unsigned( 119, 8)),3 => std_logic_vector(to_unsigned( 113, 8)),4 => std_logic_vector(to_unsigned( 100, 8)),5 => std_logic_vector(to_unsigned( 68, 8)),6 => std_logic_vector(to_unsigned( 93, 8)),7 => std_logic_vector(to_unsigned( 17, 8)),8 => std_logic_vector(to_unsigned( 107, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 442) then
				RAM <= (0 => std_logic_vector(to_unsigned( 112, 8)),1 => std_logic_vector(to_unsigned( 19, 8)),2 => std_logic_vector(to_unsigned( 44, 8)),3 => std_logic_vector(to_unsigned( 2, 8)),4 => std_logic_vector(to_unsigned( 48, 8)),5 => std_logic_vector(to_unsigned( 40, 8)),6 => std_logic_vector(to_unsigned( 14, 8)),7 => std_logic_vector(to_unsigned( 71, 8)),8 => std_logic_vector(to_unsigned( 12, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 443) then
				RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),1 => std_logic_vector(to_unsigned( 77, 8)),2 => std_logic_vector(to_unsigned( 30, 8)),3 => std_logic_vector(to_unsigned( 94, 8)),4 => std_logic_vector(to_unsigned( 54, 8)),5 => std_logic_vector(to_unsigned( 34, 8)),6 => std_logic_vector(to_unsigned( 99, 8)),7 => std_logic_vector(to_unsigned( 22, 8)),8 => std_logic_vector(to_unsigned( 59, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 444) then
				RAM <= (0 => std_logic_vector(to_unsigned( 3, 8)),1 => std_logic_vector(to_unsigned( 112, 8)),2 => std_logic_vector(to_unsigned( 20, 8)),3 => std_logic_vector(to_unsigned( 106, 8)),4 => std_logic_vector(to_unsigned( 119, 8)),5 => std_logic_vector(to_unsigned( 102, 8)),6 => std_logic_vector(to_unsigned( 65, 8)),7 => std_logic_vector(to_unsigned( 41, 8)),8 => std_logic_vector(to_unsigned( 24, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 445) then
				RAM <= (0 => std_logic_vector(to_unsigned( 1, 8)),1 => std_logic_vector(to_unsigned( 45, 8)),2 => std_logic_vector(to_unsigned( 50, 8)),3 => std_logic_vector(to_unsigned( 8, 8)),4 => std_logic_vector(to_unsigned( 75, 8)),5 => std_logic_vector(to_unsigned( 18, 8)),6 => std_logic_vector(to_unsigned( 97, 8)),7 => std_logic_vector(to_unsigned( 89, 8)),8 => std_logic_vector(to_unsigned( 42, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 446) then
				RAM <= (0 => std_logic_vector(to_unsigned( 6, 8)),1 => std_logic_vector(to_unsigned( 48, 8)),2 => std_logic_vector(to_unsigned( 40, 8)),3 => std_logic_vector(to_unsigned( 74, 8)),4 => std_logic_vector(to_unsigned( 68, 8)),5 => std_logic_vector(to_unsigned( 11, 8)),6 => std_logic_vector(to_unsigned( 30, 8)),7 => std_logic_vector(to_unsigned( 17, 8)),8 => std_logic_vector(to_unsigned( 45, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 447) then
				RAM <= (0 => std_logic_vector(to_unsigned( 31, 8)),1 => std_logic_vector(to_unsigned( 46, 8)),2 => std_logic_vector(to_unsigned( 61, 8)),3 => std_logic_vector(to_unsigned( 71, 8)),4 => std_logic_vector(to_unsigned( 8, 8)),5 => std_logic_vector(to_unsigned( 65, 8)),6 => std_logic_vector(to_unsigned( 94, 8)),7 => std_logic_vector(to_unsigned( 12, 8)),8 => std_logic_vector(to_unsigned( 50, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 448) then
				RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),1 => std_logic_vector(to_unsigned( 91, 8)),2 => std_logic_vector(to_unsigned( 73, 8)),3 => std_logic_vector(to_unsigned( 56, 8)),4 => std_logic_vector(to_unsigned( 102, 8)),5 => std_logic_vector(to_unsigned( 61, 8)),6 => std_logic_vector(to_unsigned( 85, 8)),7 => std_logic_vector(to_unsigned( 112, 8)),8 => std_logic_vector(to_unsigned( 63, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 449) then
				RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),1 => std_logic_vector(to_unsigned( 114, 8)),2 => std_logic_vector(to_unsigned( 108, 8)),3 => std_logic_vector(to_unsigned( 75, 8)),4 => std_logic_vector(to_unsigned( 23, 8)),5 => std_logic_vector(to_unsigned( 9, 8)),6 => std_logic_vector(to_unsigned( 30, 8)),7 => std_logic_vector(to_unsigned( 43, 8)),8 => std_logic_vector(to_unsigned( 79, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 450) then
				RAM <= (0 => std_logic_vector(to_unsigned( 62, 8)),1 => std_logic_vector(to_unsigned( 96, 8)),2 => std_logic_vector(to_unsigned( 32, 8)),3 => std_logic_vector(to_unsigned( 42, 8)),4 => std_logic_vector(to_unsigned( 82, 8)),5 => std_logic_vector(to_unsigned( 116, 8)),6 => std_logic_vector(to_unsigned( 78, 8)),7 => std_logic_vector(to_unsigned( 10, 8)),8 => std_logic_vector(to_unsigned( 110, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 451) then
				RAM <= (0 => std_logic_vector(to_unsigned( 18, 8)),1 => std_logic_vector(to_unsigned( 56, 8)),2 => std_logic_vector(to_unsigned( 90, 8)),3 => std_logic_vector(to_unsigned( 69, 8)),4 => std_logic_vector(to_unsigned( 124, 8)),5 => std_logic_vector(to_unsigned( 117, 8)),6 => std_logic_vector(to_unsigned( 26, 8)),7 => std_logic_vector(to_unsigned( 103, 8)),8 => std_logic_vector(to_unsigned( 78, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 452) then
				RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),1 => std_logic_vector(to_unsigned( 11, 8)),2 => std_logic_vector(to_unsigned( 80, 8)),3 => std_logic_vector(to_unsigned( 102, 8)),4 => std_logic_vector(to_unsigned( 43, 8)),5 => std_logic_vector(to_unsigned( 4, 8)),6 => std_logic_vector(to_unsigned( 69, 8)),7 => std_logic_vector(to_unsigned( 25, 8)),8 => std_logic_vector(to_unsigned( 7, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 453) then
				RAM <= (0 => std_logic_vector(to_unsigned( 10, 8)),1 => std_logic_vector(to_unsigned( 64, 8)),2 => std_logic_vector(to_unsigned( 0, 8)),3 => std_logic_vector(to_unsigned( 74, 8)),4 => std_logic_vector(to_unsigned( 78, 8)),5 => std_logic_vector(to_unsigned( 42, 8)),6 => std_logic_vector(to_unsigned( 120, 8)),7 => std_logic_vector(to_unsigned( 112, 8)),8 => std_logic_vector(to_unsigned( 121, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 454) then
				RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),1 => std_logic_vector(to_unsigned( 7, 8)),2 => std_logic_vector(to_unsigned( 2, 8)),3 => std_logic_vector(to_unsigned( 117, 8)),4 => std_logic_vector(to_unsigned( 24, 8)),5 => std_logic_vector(to_unsigned( 32, 8)),6 => std_logic_vector(to_unsigned( 44, 8)),7 => std_logic_vector(to_unsigned( 95, 8)),8 => std_logic_vector(to_unsigned( 62, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 455) then
				RAM <= (0 => std_logic_vector(to_unsigned( 105, 8)),1 => std_logic_vector(to_unsigned( 83, 8)),2 => std_logic_vector(to_unsigned( 38, 8)),3 => std_logic_vector(to_unsigned( 14, 8)),4 => std_logic_vector(to_unsigned( 110, 8)),5 => std_logic_vector(to_unsigned( 59, 8)),6 => std_logic_vector(to_unsigned( 124, 8)),7 => std_logic_vector(to_unsigned( 63, 8)),8 => std_logic_vector(to_unsigned( 18, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 456) then
				RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 46, 8)),3 => std_logic_vector(to_unsigned( 12, 8)),4 => std_logic_vector(to_unsigned( 17, 8)),5 => std_logic_vector(to_unsigned( 63, 8)),6 => std_logic_vector(to_unsigned( 73, 8)),7 => std_logic_vector(to_unsigned( 56, 8)),8 => std_logic_vector(to_unsigned( 42, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 457) then
				RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),1 => std_logic_vector(to_unsigned( 53, 8)),2 => std_logic_vector(to_unsigned( 20, 8)),3 => std_logic_vector(to_unsigned( 43, 8)),4 => std_logic_vector(to_unsigned( 24, 8)),5 => std_logic_vector(to_unsigned( 8, 8)),6 => std_logic_vector(to_unsigned( 35, 8)),7 => std_logic_vector(to_unsigned( 99, 8)),8 => std_logic_vector(to_unsigned( 85, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 458) then
				RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),1 => std_logic_vector(to_unsigned( 93, 8)),2 => std_logic_vector(to_unsigned( 83, 8)),3 => std_logic_vector(to_unsigned( 78, 8)),4 => std_logic_vector(to_unsigned( 63, 8)),5 => std_logic_vector(to_unsigned( 109, 8)),6 => std_logic_vector(to_unsigned( 74, 8)),7 => std_logic_vector(to_unsigned( 14, 8)),8 => std_logic_vector(to_unsigned( 45, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 459) then
				RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),1 => std_logic_vector(to_unsigned( 32, 8)),2 => std_logic_vector(to_unsigned( 79, 8)),3 => std_logic_vector(to_unsigned( 10, 8)),4 => std_logic_vector(to_unsigned( 74, 8)),5 => std_logic_vector(to_unsigned( 88, 8)),6 => std_logic_vector(to_unsigned( 122, 8)),7 => std_logic_vector(to_unsigned( 66, 8)),8 => std_logic_vector(to_unsigned( 111, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 460) then
				RAM <= (0 => std_logic_vector(to_unsigned( 14, 8)),1 => std_logic_vector(to_unsigned( 23, 8)),2 => std_logic_vector(to_unsigned( 110, 8)),3 => std_logic_vector(to_unsigned( 86, 8)),4 => std_logic_vector(to_unsigned( 29, 8)),5 => std_logic_vector(to_unsigned( 99, 8)),6 => std_logic_vector(to_unsigned( 52, 8)),7 => std_logic_vector(to_unsigned( 120, 8)),8 => std_logic_vector(to_unsigned( 37, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 461) then
				RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),1 => std_logic_vector(to_unsigned( 106, 8)),2 => std_logic_vector(to_unsigned( 24, 8)),3 => std_logic_vector(to_unsigned( 123, 8)),4 => std_logic_vector(to_unsigned( 17, 8)),5 => std_logic_vector(to_unsigned( 112, 8)),6 => std_logic_vector(to_unsigned( 80, 8)),7 => std_logic_vector(to_unsigned( 8, 8)),8 => std_logic_vector(to_unsigned( 67, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 462) then
				RAM <= (0 => std_logic_vector(to_unsigned( 70, 8)),1 => std_logic_vector(to_unsigned( 115, 8)),2 => std_logic_vector(to_unsigned( 32, 8)),3 => std_logic_vector(to_unsigned( 101, 8)),4 => std_logic_vector(to_unsigned( 21, 8)),5 => std_logic_vector(to_unsigned( 107, 8)),6 => std_logic_vector(to_unsigned( 111, 8)),7 => std_logic_vector(to_unsigned( 7, 8)),8 => std_logic_vector(to_unsigned( 19, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 463) then
				RAM <= (0 => std_logic_vector(to_unsigned( 73, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 82, 8)),3 => std_logic_vector(to_unsigned( 21, 8)),4 => std_logic_vector(to_unsigned( 109, 8)),5 => std_logic_vector(to_unsigned( 0, 8)),6 => std_logic_vector(to_unsigned( 41, 8)),7 => std_logic_vector(to_unsigned( 89, 8)),8 => std_logic_vector(to_unsigned( 59, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 464) then
				RAM <= (0 => std_logic_vector(to_unsigned( 63, 8)),1 => std_logic_vector(to_unsigned( 58, 8)),2 => std_logic_vector(to_unsigned( 111, 8)),3 => std_logic_vector(to_unsigned( 99, 8)),4 => std_logic_vector(to_unsigned( 9, 8)),5 => std_logic_vector(to_unsigned( 85, 8)),6 => std_logic_vector(to_unsigned( 93, 8)),7 => std_logic_vector(to_unsigned( 106, 8)),8 => std_logic_vector(to_unsigned( 113, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 465) then
				RAM <= (0 => std_logic_vector(to_unsigned( 2, 8)),1 => std_logic_vector(to_unsigned( 26, 8)),2 => std_logic_vector(to_unsigned( 77, 8)),3 => std_logic_vector(to_unsigned( 124, 8)),4 => std_logic_vector(to_unsigned( 61, 8)),5 => std_logic_vector(to_unsigned( 11, 8)),6 => std_logic_vector(to_unsigned( 50, 8)),7 => std_logic_vector(to_unsigned( 22, 8)),8 => std_logic_vector(to_unsigned( 94, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 466) then
				RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),1 => std_logic_vector(to_unsigned( 85, 8)),2 => std_logic_vector(to_unsigned( 20, 8)),3 => std_logic_vector(to_unsigned( 0, 8)),4 => std_logic_vector(to_unsigned( 9, 8)),5 => std_logic_vector(to_unsigned( 99, 8)),6 => std_logic_vector(to_unsigned( 63, 8)),7 => std_logic_vector(to_unsigned( 104, 8)),8 => std_logic_vector(to_unsigned( 30, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 467) then
				RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),1 => std_logic_vector(to_unsigned( 105, 8)),2 => std_logic_vector(to_unsigned( 1, 8)),3 => std_logic_vector(to_unsigned( 29, 8)),4 => std_logic_vector(to_unsigned( 110, 8)),5 => std_logic_vector(to_unsigned( 66, 8)),6 => std_logic_vector(to_unsigned( 43, 8)),7 => std_logic_vector(to_unsigned( 12, 8)),8 => std_logic_vector(to_unsigned( 39, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 468) then
				RAM <= (0 => std_logic_vector(to_unsigned( 116, 8)),1 => std_logic_vector(to_unsigned( 95, 8)),2 => std_logic_vector(to_unsigned( 11, 8)),3 => std_logic_vector(to_unsigned( 105, 8)),4 => std_logic_vector(to_unsigned( 48, 8)),5 => std_logic_vector(to_unsigned( 77, 8)),6 => std_logic_vector(to_unsigned( 63, 8)),7 => std_logic_vector(to_unsigned( 32, 8)),8 => std_logic_vector(to_unsigned( 5, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 469) then
				RAM <= (0 => std_logic_vector(to_unsigned( 108, 8)),1 => std_logic_vector(to_unsigned( 98, 8)),2 => std_logic_vector(to_unsigned( 30, 8)),3 => std_logic_vector(to_unsigned( 51, 8)),4 => std_logic_vector(to_unsigned( 10, 8)),5 => std_logic_vector(to_unsigned( 121, 8)),6 => std_logic_vector(to_unsigned( 21, 8)),7 => std_logic_vector(to_unsigned( 73, 8)),8 => std_logic_vector(to_unsigned( 65, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 470) then
				RAM <= (0 => std_logic_vector(to_unsigned( 64, 8)),1 => std_logic_vector(to_unsigned( 59, 8)),2 => std_logic_vector(to_unsigned( 75, 8)),3 => std_logic_vector(to_unsigned( 118, 8)),4 => std_logic_vector(to_unsigned( 91, 8)),5 => std_logic_vector(to_unsigned( 111, 8)),6 => std_logic_vector(to_unsigned( 3, 8)),7 => std_logic_vector(to_unsigned( 8, 8)),8 => std_logic_vector(to_unsigned( 6, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 471) then
				RAM <= (0 => std_logic_vector(to_unsigned( 113, 8)),1 => std_logic_vector(to_unsigned( 10, 8)),2 => std_logic_vector(to_unsigned( 50, 8)),3 => std_logic_vector(to_unsigned( 23, 8)),4 => std_logic_vector(to_unsigned( 14, 8)),5 => std_logic_vector(to_unsigned( 43, 8)),6 => std_logic_vector(to_unsigned( 85, 8)),7 => std_logic_vector(to_unsigned( 108, 8)),8 => std_logic_vector(to_unsigned( 95, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 472) then
				RAM <= (0 => std_logic_vector(to_unsigned( 118, 8)),1 => std_logic_vector(to_unsigned( 63, 8)),2 => std_logic_vector(to_unsigned( 76, 8)),3 => std_logic_vector(to_unsigned( 23, 8)),4 => std_logic_vector(to_unsigned( 32, 8)),5 => std_logic_vector(to_unsigned( 99, 8)),6 => std_logic_vector(to_unsigned( 45, 8)),7 => std_logic_vector(to_unsigned( 5, 8)),8 => std_logic_vector(to_unsigned( 105, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 473) then
				RAM <= (0 => std_logic_vector(to_unsigned( 111, 8)),1 => std_logic_vector(to_unsigned( 55, 8)),2 => std_logic_vector(to_unsigned( 105, 8)),3 => std_logic_vector(to_unsigned( 119, 8)),4 => std_logic_vector(to_unsigned( 7, 8)),5 => std_logic_vector(to_unsigned( 95, 8)),6 => std_logic_vector(to_unsigned( 18, 8)),7 => std_logic_vector(to_unsigned( 80, 8)),8 => std_logic_vector(to_unsigned( 40, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 474) then
				RAM <= (0 => std_logic_vector(to_unsigned( 58, 8)),1 => std_logic_vector(to_unsigned( 53, 8)),2 => std_logic_vector(to_unsigned( 102, 8)),3 => std_logic_vector(to_unsigned( 71, 8)),4 => std_logic_vector(to_unsigned( 8, 8)),5 => std_logic_vector(to_unsigned( 28, 8)),6 => std_logic_vector(to_unsigned( 16, 8)),7 => std_logic_vector(to_unsigned( 121, 8)),8 => std_logic_vector(to_unsigned( 93, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 475) then
				RAM <= (0 => std_logic_vector(to_unsigned( 70, 8)),1 => std_logic_vector(to_unsigned( 62, 8)),2 => std_logic_vector(to_unsigned( 98, 8)),3 => std_logic_vector(to_unsigned( 53, 8)),4 => std_logic_vector(to_unsigned( 26, 8)),5 => std_logic_vector(to_unsigned( 9, 8)),6 => std_logic_vector(to_unsigned( 102, 8)),7 => std_logic_vector(to_unsigned( 88, 8)),8 => std_logic_vector(to_unsigned( 61, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 476) then
				RAM <= (0 => std_logic_vector(to_unsigned( 112, 8)),1 => std_logic_vector(to_unsigned( 25, 8)),2 => std_logic_vector(to_unsigned( 59, 8)),3 => std_logic_vector(to_unsigned( 54, 8)),4 => std_logic_vector(to_unsigned( 43, 8)),5 => std_logic_vector(to_unsigned( 31, 8)),6 => std_logic_vector(to_unsigned( 117, 8)),7 => std_logic_vector(to_unsigned( 65, 8)),8 => std_logic_vector(to_unsigned( 57, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 477) then
				RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),1 => std_logic_vector(to_unsigned( 69, 8)),2 => std_logic_vector(to_unsigned( 86, 8)),3 => std_logic_vector(to_unsigned( 51, 8)),4 => std_logic_vector(to_unsigned( 41, 8)),5 => std_logic_vector(to_unsigned( 22, 8)),6 => std_logic_vector(to_unsigned( 90, 8)),7 => std_logic_vector(to_unsigned( 113, 8)),8 => std_logic_vector(to_unsigned( 28, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 478) then
				RAM <= (0 => std_logic_vector(to_unsigned( 106, 8)),1 => std_logic_vector(to_unsigned( 27, 8)),2 => std_logic_vector(to_unsigned( 18, 8)),3 => std_logic_vector(to_unsigned( 123, 8)),4 => std_logic_vector(to_unsigned( 82, 8)),5 => std_logic_vector(to_unsigned( 44, 8)),6 => std_logic_vector(to_unsigned( 3, 8)),7 => std_logic_vector(to_unsigned( 94, 8)),8 => std_logic_vector(to_unsigned( 29, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 479) then
				RAM <= (0 => std_logic_vector(to_unsigned( 23, 8)),1 => std_logic_vector(to_unsigned( 120, 8)),2 => std_logic_vector(to_unsigned( 100, 8)),3 => std_logic_vector(to_unsigned( 83, 8)),4 => std_logic_vector(to_unsigned( 110, 8)),5 => std_logic_vector(to_unsigned( 48, 8)),6 => std_logic_vector(to_unsigned( 94, 8)),7 => std_logic_vector(to_unsigned( 13, 8)),8 => std_logic_vector(to_unsigned( 7, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 480) then
				RAM <= (0 => std_logic_vector(to_unsigned( 120, 8)),1 => std_logic_vector(to_unsigned( 91, 8)),2 => std_logic_vector(to_unsigned( 57, 8)),3 => std_logic_vector(to_unsigned( 40, 8)),4 => std_logic_vector(to_unsigned( 6, 8)),5 => std_logic_vector(to_unsigned( 124, 8)),6 => std_logic_vector(to_unsigned( 80, 8)),7 => std_logic_vector(to_unsigned( 34, 8)),8 => std_logic_vector(to_unsigned( 127, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 481) then
				RAM <= (0 => std_logic_vector(to_unsigned( 75, 8)),1 => std_logic_vector(to_unsigned( 5, 8)),2 => std_logic_vector(to_unsigned( 24, 8)),3 => std_logic_vector(to_unsigned( 107, 8)),4 => std_logic_vector(to_unsigned( 71, 8)),5 => std_logic_vector(to_unsigned( 50, 8)),6 => std_logic_vector(to_unsigned( 82, 8)),7 => std_logic_vector(to_unsigned( 30, 8)),8 => std_logic_vector(to_unsigned( 24, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 482) then
				RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),1 => std_logic_vector(to_unsigned( 8, 8)),2 => std_logic_vector(to_unsigned( 112, 8)),3 => std_logic_vector(to_unsigned( 65, 8)),4 => std_logic_vector(to_unsigned( 119, 8)),5 => std_logic_vector(to_unsigned( 27, 8)),6 => std_logic_vector(to_unsigned( 3, 8)),7 => std_logic_vector(to_unsigned( 107, 8)),8 => std_logic_vector(to_unsigned( 125, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 483) then
				RAM <= (0 => std_logic_vector(to_unsigned( 93, 8)),1 => std_logic_vector(to_unsigned( 15, 8)),2 => std_logic_vector(to_unsigned( 19, 8)),3 => std_logic_vector(to_unsigned( 114, 8)),4 => std_logic_vector(to_unsigned( 78, 8)),5 => std_logic_vector(to_unsigned( 8, 8)),6 => std_logic_vector(to_unsigned( 85, 8)),7 => std_logic_vector(to_unsigned( 36, 8)),8 => std_logic_vector(to_unsigned( 85, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 484) then
				RAM <= (0 => std_logic_vector(to_unsigned( 50, 8)),1 => std_logic_vector(to_unsigned( 73, 8)),2 => std_logic_vector(to_unsigned( 117, 8)),3 => std_logic_vector(to_unsigned( 1, 8)),4 => std_logic_vector(to_unsigned( 110, 8)),5 => std_logic_vector(to_unsigned( 105, 8)),6 => std_logic_vector(to_unsigned( 11, 8)),7 => std_logic_vector(to_unsigned( 92, 8)),8 => std_logic_vector(to_unsigned( 8, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 485) then
				RAM <= (0 => std_logic_vector(to_unsigned( 67, 8)),1 => std_logic_vector(to_unsigned( 75, 8)),2 => std_logic_vector(to_unsigned( 3, 8)),3 => std_logic_vector(to_unsigned( 42, 8)),4 => std_logic_vector(to_unsigned( 50, 8)),5 => std_logic_vector(to_unsigned( 15, 8)),6 => std_logic_vector(to_unsigned( 34, 8)),7 => std_logic_vector(to_unsigned( 96, 8)),8 => std_logic_vector(to_unsigned( 61, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 486) then
				RAM <= (0 => std_logic_vector(to_unsigned( 17, 8)),1 => std_logic_vector(to_unsigned( 117, 8)),2 => std_logic_vector(to_unsigned( 92, 8)),3 => std_logic_vector(to_unsigned( 8, 8)),4 => std_logic_vector(to_unsigned( 123, 8)),5 => std_logic_vector(to_unsigned( 51, 8)),6 => std_logic_vector(to_unsigned( 60, 8)),7 => std_logic_vector(to_unsigned( 73, 8)),8 => std_logic_vector(to_unsigned( 106, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 487) then
				RAM <= (0 => std_logic_vector(to_unsigned( 48, 8)),1 => std_logic_vector(to_unsigned( 3, 8)),2 => std_logic_vector(to_unsigned( 23, 8)),3 => std_logic_vector(to_unsigned( 82, 8)),4 => std_logic_vector(to_unsigned( 36, 8)),5 => std_logic_vector(to_unsigned( 61, 8)),6 => std_logic_vector(to_unsigned( 95, 8)),7 => std_logic_vector(to_unsigned( 77, 8)),8 => std_logic_vector(to_unsigned( 93, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 488) then
				RAM <= (0 => std_logic_vector(to_unsigned( 114, 8)),1 => std_logic_vector(to_unsigned( 75, 8)),2 => std_logic_vector(to_unsigned( 14, 8)),3 => std_logic_vector(to_unsigned( 93, 8)),4 => std_logic_vector(to_unsigned( 123, 8)),5 => std_logic_vector(to_unsigned( 97, 8)),6 => std_logic_vector(to_unsigned( 28, 8)),7 => std_logic_vector(to_unsigned( 55, 8)),8 => std_logic_vector(to_unsigned( 58, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 489) then
				RAM <= (0 => std_logic_vector(to_unsigned( 69, 8)),1 => std_logic_vector(to_unsigned( 48, 8)),2 => std_logic_vector(to_unsigned( 83, 8)),3 => std_logic_vector(to_unsigned( 63, 8)),4 => std_logic_vector(to_unsigned( 116, 8)),5 => std_logic_vector(to_unsigned( 53, 8)),6 => std_logic_vector(to_unsigned( 89, 8)),7 => std_logic_vector(to_unsigned( 106, 8)),8 => std_logic_vector(to_unsigned( 57, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 490) then
				RAM <= (0 => std_logic_vector(to_unsigned( 32, 8)),1 => std_logic_vector(to_unsigned( 105, 8)),2 => std_logic_vector(to_unsigned( 44, 8)),3 => std_logic_vector(to_unsigned( 21, 8)),4 => std_logic_vector(to_unsigned( 12, 8)),5 => std_logic_vector(to_unsigned( 110, 8)),6 => std_logic_vector(to_unsigned( 70, 8)),7 => std_logic_vector(to_unsigned( 39, 8)),8 => std_logic_vector(to_unsigned( 12, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 491) then
				RAM <= (0 => std_logic_vector(to_unsigned( 81, 8)),1 => std_logic_vector(to_unsigned( 53, 8)),2 => std_logic_vector(to_unsigned( 16, 8)),3 => std_logic_vector(to_unsigned( 33, 8)),4 => std_logic_vector(to_unsigned( 107, 8)),5 => std_logic_vector(to_unsigned( 4, 8)),6 => std_logic_vector(to_unsigned( 60, 8)),7 => std_logic_vector(to_unsigned( 88, 8)),8 => std_logic_vector(to_unsigned( 26, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 492) then
				RAM <= (0 => std_logic_vector(to_unsigned( 0, 8)),1 => std_logic_vector(to_unsigned( 6, 8)),2 => std_logic_vector(to_unsigned( 18, 8)),3 => std_logic_vector(to_unsigned( 82, 8)),4 => std_logic_vector(to_unsigned( 115, 8)),5 => std_logic_vector(to_unsigned( 124, 8)),6 => std_logic_vector(to_unsigned( 51, 8)),7 => std_logic_vector(to_unsigned( 107, 8)),8 => std_logic_vector(to_unsigned( 1, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 493) then
				RAM <= (0 => std_logic_vector(to_unsigned( 59, 8)),1 => std_logic_vector(to_unsigned( 88, 8)),2 => std_logic_vector(to_unsigned( 55, 8)),3 => std_logic_vector(to_unsigned( 123, 8)),4 => std_logic_vector(to_unsigned( 116, 8)),5 => std_logic_vector(to_unsigned( 21, 8)),6 => std_logic_vector(to_unsigned( 44, 8)),7 => std_logic_vector(to_unsigned( 78, 8)),8 => std_logic_vector(to_unsigned( 125, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 494) then
				RAM <= (0 => std_logic_vector(to_unsigned( 66, 8)),1 => std_logic_vector(to_unsigned( 74, 8)),2 => std_logic_vector(to_unsigned( 93, 8)),3 => std_logic_vector(to_unsigned( 98, 8)),4 => std_logic_vector(to_unsigned( 31, 8)),5 => std_logic_vector(to_unsigned( 6, 8)),6 => std_logic_vector(to_unsigned( 83, 8)),7 => std_logic_vector(to_unsigned( 61, 8)),8 => std_logic_vector(to_unsigned( 52, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 495) then
				RAM <= (0 => std_logic_vector(to_unsigned( 37, 8)),1 => std_logic_vector(to_unsigned( 101, 8)),2 => std_logic_vector(to_unsigned( 44, 8)),3 => std_logic_vector(to_unsigned( 23, 8)),4 => std_logic_vector(to_unsigned( 118, 8)),5 => std_logic_vector(to_unsigned( 65, 8)),6 => std_logic_vector(to_unsigned( 28, 8)),7 => std_logic_vector(to_unsigned( 85, 8)),8 => std_logic_vector(to_unsigned( 126, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 496) then
				RAM <= (0 => std_logic_vector(to_unsigned( 124, 8)),1 => std_logic_vector(to_unsigned( 50, 8)),2 => std_logic_vector(to_unsigned( 24, 8)),3 => std_logic_vector(to_unsigned( 91, 8)),4 => std_logic_vector(to_unsigned( 5, 8)),5 => std_logic_vector(to_unsigned( 108, 8)),6 => std_logic_vector(to_unsigned( 11, 8)),7 => std_logic_vector(to_unsigned( 44, 8)),8 => std_logic_vector(to_unsigned( 36, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 497) then
				RAM <= (0 => std_logic_vector(to_unsigned( 122, 8)),1 => std_logic_vector(to_unsigned( 100, 8)),2 => std_logic_vector(to_unsigned( 21, 8)),3 => std_logic_vector(to_unsigned( 6, 8)),4 => std_logic_vector(to_unsigned( 78, 8)),5 => std_logic_vector(to_unsigned( 25, 8)),6 => std_logic_vector(to_unsigned( 56, 8)),7 => std_logic_vector(to_unsigned( 0, 8)),8 => std_logic_vector(to_unsigned( 52, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			elsif(numero_test = 498) then
				RAM <= (0 => std_logic_vector(to_unsigned( 82, 8)),1 => std_logic_vector(to_unsigned( 100, 8)),2 => std_logic_vector(to_unsigned( 13, 8)),3 => std_logic_vector(to_unsigned( 25, 8)),4 => std_logic_vector(to_unsigned( 88, 8)),5 => std_logic_vector(to_unsigned( 34, 8)),6 => std_logic_vector(to_unsigned( 59, 8)),7 => std_logic_vector(to_unsigned( 53, 8)),8 => std_logic_vector(to_unsigned( 90, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			else
				RAM <= (0 => std_logic_vector(to_unsigned( 44, 8)),1 => std_logic_vector(to_unsigned( 11, 8)),2 => std_logic_vector(to_unsigned( 36, 8)),3 => std_logic_vector(to_unsigned( 95, 8)),4 => std_logic_vector(to_unsigned( 3, 8)),5 => std_logic_vector(to_unsigned( 121, 8)),6 => std_logic_vector(to_unsigned( 113, 8)),7 => std_logic_vector(to_unsigned( 102, 8)),8 => std_logic_vector(to_unsigned( 106, 8)), others => (others =>'0'));
				numero_test := numero_test+1;
			end if;
		end if;
	end if;
end process;


test : process is

	begin

		-- test numero 0

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(32 , 8)) report "TEST FALLITO. Expected  32  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 0 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 1

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(129 , 8)) report "TEST FALLITO. Expected  129  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 1 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 2

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(75 , 8)) report "TEST FALLITO. Expected  75  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 2 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 3

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(248 , 8)) report "TEST FALLITO. Expected  248  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 3 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 4

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(118 , 8)) report "TEST FALLITO. Expected  118  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 4 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 5

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(35 , 8)) report "TEST FALLITO. Expected  35  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 5 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 6

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(180 , 8)) report "TEST FALLITO. Expected  180  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 6 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 7

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(100 , 8)) report "TEST FALLITO. Expected  100  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 7 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 8

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(52 , 8)) report "TEST FALLITO. Expected  52  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 8 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 9

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(4 , 8)) report "TEST FALLITO. Expected  4  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 9 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 10

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(100 , 8)) report "TEST FALLITO. Expected  100  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 10 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 11

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(79 , 8)) report "TEST FALLITO. Expected  79  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 11 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 12

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(47 , 8)) report "TEST FALLITO. Expected  47  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 12 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 13

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(248 , 8)) report "TEST FALLITO. Expected  248  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 13 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 14

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(62 , 8)) report "TEST FALLITO. Expected  62  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 14 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 15

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(93 , 8)) report "TEST FALLITO. Expected  93  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 15 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 16

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(26 , 8)) report "TEST FALLITO. Expected  26  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 16 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 17

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(161 , 8)) report "TEST FALLITO. Expected  161  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 17 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 18

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(177 , 8)) report "TEST FALLITO. Expected  177  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 18 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 19

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(25 , 8)) report "TEST FALLITO. Expected  25  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 19 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 20

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(226 , 8)) report "TEST FALLITO. Expected  226  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 20 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 21

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(110 , 8)) report "TEST FALLITO. Expected  110  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 21 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 22

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(136 , 8)) report "TEST FALLITO. Expected  136  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 22 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 23

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(62 , 8)) report "TEST FALLITO. Expected  62  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 23 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 24

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(115 , 8)) report "TEST FALLITO. Expected  115  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 24 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 25

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(34 , 8)) report "TEST FALLITO. Expected  34  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 25 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 26

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(193 , 8)) report "TEST FALLITO. Expected  193  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 26 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 27

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(14 , 8)) report "TEST FALLITO. Expected  14  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 27 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 28

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(129 , 8)) report "TEST FALLITO. Expected  129  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 28 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 29

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(248 , 8)) report "TEST FALLITO. Expected  248  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 29 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 30

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(102 , 8)) report "TEST FALLITO. Expected  102  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 30 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 31

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(64 , 8)) report "TEST FALLITO. Expected  64  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 31 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 32

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(53 , 8)) report "TEST FALLITO. Expected  53  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 32 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 33

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(89 , 8)) report "TEST FALLITO. Expected  89  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 33 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 34

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(112 , 8)) report "TEST FALLITO. Expected  112  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 34 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 35

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(129 , 8)) report "TEST FALLITO. Expected  129  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 35 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 36

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(67 , 8)) report "TEST FALLITO. Expected  67  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 36 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 37

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(106 , 8)) report "TEST FALLITO. Expected  106  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 37 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 38

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(241 , 8)) report "TEST FALLITO. Expected  241  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 38 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 39

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(107 , 8)) report "TEST FALLITO. Expected  107  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 39 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 40

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(46 , 8)) report "TEST FALLITO. Expected  46  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 40 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 41

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(35 , 8)) report "TEST FALLITO. Expected  35  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 41 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 42

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(56 , 8)) report "TEST FALLITO. Expected  56  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 42 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 43

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(41 , 8)) report "TEST FALLITO. Expected  41  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 43 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 44

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(23 , 8)) report "TEST FALLITO. Expected  23  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 44 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 45

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(242 , 8)) report "TEST FALLITO. Expected  242  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 45 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 46

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(148 , 8)) report "TEST FALLITO. Expected  148  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 46 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 47

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(164 , 8)) report "TEST FALLITO. Expected  164  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 47 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 48 interrotto

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		--interruzione
		--wait for c_CLOCK_PERIOD;
		--wait until tb_done = '1';
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;


		-- test numero 49 asincrono

		wait for 100 ns;
		--wait for c_CLOCK_PERIOD;--------------------------il reset non arriva sul clock
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		--tb_start <= '1';----------------------------------lo start � ancora alto dal test precedente
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(116 , 8)) report "TEST FALLITO. Expected  116  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 49 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 50

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(164 , 8)) report "TEST FALLITO. Expected  164  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 50 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 51

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(72 , 8)) report "TEST FALLITO. Expected  72  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 51 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 52

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(178 , 8)) report "TEST FALLITO. Expected  178  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 52 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 53

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(244 , 8)) report "TEST FALLITO. Expected  244  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 53 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 54

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(225 , 8)) report "TEST FALLITO. Expected  225  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 54 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 55

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(59 , 8)) report "TEST FALLITO. Expected  59  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 55 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 56

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(99 , 8)) report "TEST FALLITO. Expected  99  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 56 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 57

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(94 , 8)) report "TEST FALLITO. Expected  94  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 57 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 58

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(124 , 8)) report "TEST FALLITO. Expected  124  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 58 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 59

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(31 , 8)) report "TEST FALLITO. Expected  31  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 59 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 60

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(52 , 8)) report "TEST FALLITO. Expected  52  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 60 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 61

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(44 , 8)) report "TEST FALLITO. Expected  44  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 61 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 62

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(90 , 8)) report "TEST FALLITO. Expected  90  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 62 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 63

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(0 , 8)) report "TEST FALLITO. Expected  0  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 63 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 64

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(25 , 8)) report "TEST FALLITO. Expected  25  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 64 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 65

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(115 , 8)) report "TEST FALLITO. Expected  115  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 65 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 66

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(62 , 8)) report "TEST FALLITO. Expected  62  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 66 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 67

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(4 , 8)) report "TEST FALLITO. Expected  4  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 67 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 68

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(29 , 8)) report "TEST FALLITO. Expected  29  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 68 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 69

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(82 , 8)) report "TEST FALLITO. Expected  82  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 69 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 70

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(125 , 8)) report "TEST FALLITO. Expected  125  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 70 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 71

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(162 , 8)) report "TEST FALLITO. Expected  162  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 71 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 72

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(7 , 8)) report "TEST FALLITO. Expected  7  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 72 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 73

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(37 , 8)) report "TEST FALLITO. Expected  37  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 73 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 74

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(69 , 8)) report "TEST FALLITO. Expected  69  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 74 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 75

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(18 , 8)) report "TEST FALLITO. Expected  18  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 75 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 76

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(88 , 8)) report "TEST FALLITO. Expected  88  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 76 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 77

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(58 , 8)) report "TEST FALLITO. Expected  58  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 77 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 78

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(177 , 8)) report "TEST FALLITO. Expected  177  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 78 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 79

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(112 , 8)) report "TEST FALLITO. Expected  112  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 79 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 80

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(27 , 8)) report "TEST FALLITO. Expected  27  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 80 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 81

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(24 , 8)) report "TEST FALLITO. Expected  24  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 81 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 82

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(90 , 8)) report "TEST FALLITO. Expected  90  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 82 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 83

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(130 , 8)) report "TEST FALLITO. Expected  130  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 83 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 84

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(209 , 8)) report "TEST FALLITO. Expected  209  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 84 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 85

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(226 , 8)) report "TEST FALLITO. Expected  226  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 85 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 86

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(31 , 8)) report "TEST FALLITO. Expected  31  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 86 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 87

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(121 , 8)) report "TEST FALLITO. Expected  121  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 87 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 88

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(60 , 8)) report "TEST FALLITO. Expected  60  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 88 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 89

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(242 , 8)) report "TEST FALLITO. Expected  242  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 89 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 90

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(112 , 8)) report "TEST FALLITO. Expected  112  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 90 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 91

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(68 , 8)) report "TEST FALLITO. Expected  68  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 91 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 92

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(99 , 8)) report "TEST FALLITO. Expected  99  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 92 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 93

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(37 , 8)) report "TEST FALLITO. Expected  37  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 93 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 94

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(27 , 8)) report "TEST FALLITO. Expected  27  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 94 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 95

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(30 , 8)) report "TEST FALLITO. Expected  30  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 95 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 96

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(50 , 8)) report "TEST FALLITO. Expected  50  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 96 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 97

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(82 , 8)) report "TEST FALLITO. Expected  82  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 97 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 98 interrotto

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		--test interrotto prima di uno start
		
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '1';
		--wait for c_CLOCK_PERIOD;
		--wait until tb_done = '1';
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(161 , 8)) report "TEST FALLITO. Expected  161  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 98 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 99 asincrono

		wait for 100 ns;
		--wait for c_CLOCK_PERIOD;---------------il reset non arriva sul clock
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(77 , 8)) report "TEST FALLITO. Expected  77  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 99 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 100

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(2 , 8)) report "TEST FALLITO. Expected  2  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 100 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 101

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(19 , 8)) report "TEST FALLITO. Expected  19  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 101 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 102

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(209 , 8)) report "TEST FALLITO. Expected  209  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 102 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 103

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(72 , 8)) report "TEST FALLITO. Expected  72  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 103 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 104

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(136 , 8)) report "TEST FALLITO. Expected  136  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 104 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 105

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(58 , 8)) report "TEST FALLITO. Expected  58  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 105 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 106

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(109 , 8)) report "TEST FALLITO. Expected  109  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 106 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 107

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(168 , 8)) report "TEST FALLITO. Expected  168  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 107 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 108

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(7 , 8)) report "TEST FALLITO. Expected  7  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 108 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 109

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(89 , 8)) report "TEST FALLITO. Expected  89  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 109 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 110

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(162 , 8)) report "TEST FALLITO. Expected  162  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 110 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 111

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(88 , 8)) report "TEST FALLITO. Expected  88  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 111 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 112

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(226 , 8)) report "TEST FALLITO. Expected  226  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 112 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 113

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(11 , 8)) report "TEST FALLITO. Expected  11  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 113 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 114

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(55 , 8)) report "TEST FALLITO. Expected  55  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 114 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 115

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(10 , 8)) report "TEST FALLITO. Expected  10  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 115 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 116

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(3 , 8)) report "TEST FALLITO. Expected  3  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 116 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 117

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(57 , 8)) report "TEST FALLITO. Expected  57  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 117 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 118

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(64 , 8)) report "TEST FALLITO. Expected  64  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 118 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 119

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(13 , 8)) report "TEST FALLITO. Expected  13  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 119 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 120

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(27 , 8)) report "TEST FALLITO. Expected  27  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 120 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 121

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(74 , 8)) report "TEST FALLITO. Expected  74  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 121 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 122

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(193 , 8)) report "TEST FALLITO. Expected  193  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 122 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 123

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(72 , 8)) report "TEST FALLITO. Expected  72  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 123 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 124

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(83 , 8)) report "TEST FALLITO. Expected  83  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 124 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 125

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(226 , 8)) report "TEST FALLITO. Expected  226  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 125 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 126

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(48 , 8)) report "TEST FALLITO. Expected  48  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 126 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 127

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(41 , 8)) report "TEST FALLITO. Expected  41  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 127 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 128

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(17 , 8)) report "TEST FALLITO. Expected  17  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 128 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 129

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(216 , 8)) report "TEST FALLITO. Expected  216  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 129 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 130

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(132 , 8)) report "TEST FALLITO. Expected  132  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 130 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 131

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(93 , 8)) report "TEST FALLITO. Expected  93  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 131 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 132

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(17 , 8)) report "TEST FALLITO. Expected  17  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 132 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 133

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(41 , 8)) report "TEST FALLITO. Expected  41  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 133 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 134

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(161 , 8)) report "TEST FALLITO. Expected  161  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 134 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 135

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(40 , 8)) report "TEST FALLITO. Expected  40  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 135 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 136

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(23 , 8)) report "TEST FALLITO. Expected  23  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 136 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 137

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(31 , 8)) report "TEST FALLITO. Expected  31  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 137 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 138

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(96 , 8)) report "TEST FALLITO. Expected  96  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 138 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 139

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(3 , 8)) report "TEST FALLITO. Expected  3  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 139 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 140

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(209 , 8)) report "TEST FALLITO. Expected  209  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 140 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 141

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(112 , 8)) report "TEST FALLITO. Expected  112  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 141 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 142

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(132 , 8)) report "TEST FALLITO. Expected  132  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 142 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 143

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(132 , 8)) report "TEST FALLITO. Expected  132  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 143 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 144

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(25 , 8)) report "TEST FALLITO. Expected  25  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 144 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 145

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(40 , 8)) report "TEST FALLITO. Expected  40  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 145 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 146

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(56 , 8)) report "TEST FALLITO. Expected  56  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 146 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 147

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(56 , 8)) report "TEST FALLITO. Expected  56  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 147 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 148 interrotto

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		--interruzione specificamente dopo che � stato alzato o_done
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(58 , 8)) report "TEST FALLITO. Expected  58  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 148 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 149 asincrono

		wait for 10 ns;-------------------------attesa breve
		--wait for c_CLOCK_PERIOD;--------------reset non arriva sul clock
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(209 , 8)) report "TEST FALLITO. Expected  209  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 149 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 150

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(47 , 8)) report "TEST FALLITO. Expected  47  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 150 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 151

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(11 , 8)) report "TEST FALLITO. Expected  11  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 151 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 152

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(21 , 8)) report "TEST FALLITO. Expected  21  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 152 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 153

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(10 , 8)) report "TEST FALLITO. Expected  10  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 153 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 154

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(56 , 8)) report "TEST FALLITO. Expected  56  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 154 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 155

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(49 , 8)) report "TEST FALLITO. Expected  49  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 155 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 156

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(17 , 8)) report "TEST FALLITO. Expected  17  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 156 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 157

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(41 , 8)) report "TEST FALLITO. Expected  41  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 157 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 158

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(2 , 8)) report "TEST FALLITO. Expected  2  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 158 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 159

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(61 , 8)) report "TEST FALLITO. Expected  61  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 159 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 160

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(71 , 8)) report "TEST FALLITO. Expected  71  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 160 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 161

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(126 , 8)) report "TEST FALLITO. Expected  126  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 161 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 162

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(33 , 8)) report "TEST FALLITO. Expected  33  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 162 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 163

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(39 , 8)) report "TEST FALLITO. Expected  39  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 163 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 164

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(194 , 8)) report "TEST FALLITO. Expected  194  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 164 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 165

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(101 , 8)) report "TEST FALLITO. Expected  101  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 165 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 166

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(95 , 8)) report "TEST FALLITO. Expected  95  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 166 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 167

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(196 , 8)) report "TEST FALLITO. Expected  196  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 167 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 168

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(36 , 8)) report "TEST FALLITO. Expected  36  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 168 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 169

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(44 , 8)) report "TEST FALLITO. Expected  44  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 169 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 170

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(77 , 8)) report "TEST FALLITO. Expected  77  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 170 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 171

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(64 , 8)) report "TEST FALLITO. Expected  64  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 171 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 172

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(146 , 8)) report "TEST FALLITO. Expected  146  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 172 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 173

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(90 , 8)) report "TEST FALLITO. Expected  90  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 173 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 174

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(226 , 8)) report "TEST FALLITO. Expected  226  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 174 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 175

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(97 , 8)) report "TEST FALLITO. Expected  97  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 175 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 176

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(70 , 8)) report "TEST FALLITO. Expected  70  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 176 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 177

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(107 , 8)) report "TEST FALLITO. Expected  107  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 177 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 178

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(64 , 8)) report "TEST FALLITO. Expected  64  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 178 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 179

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(47 , 8)) report "TEST FALLITO. Expected  47  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 179 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 180

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(84 , 8)) report "TEST FALLITO. Expected  84  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 180 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 181

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(145 , 8)) report "TEST FALLITO. Expected  145  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 181 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 182

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(10 , 8)) report "TEST FALLITO. Expected  10  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 182 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 183

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(92 , 8)) report "TEST FALLITO. Expected  92  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 183 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 184

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(129 , 8)) report "TEST FALLITO. Expected  129  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 184 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 185

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(66 , 8)) report "TEST FALLITO. Expected  66  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 185 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 186

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(132 , 8)) report "TEST FALLITO. Expected  132  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 186 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 187

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(26 , 8)) report "TEST FALLITO. Expected  26  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 187 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 188

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(118 , 8)) report "TEST FALLITO. Expected  118  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 188 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 189

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(87 , 8)) report "TEST FALLITO. Expected  87  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 189 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 190

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(67 , 8)) report "TEST FALLITO. Expected  67  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 190 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 191

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(145 , 8)) report "TEST FALLITO. Expected  145  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 191 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 192

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(108 , 8)) report "TEST FALLITO. Expected  108  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 192 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 193

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(148 , 8)) report "TEST FALLITO. Expected  148  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 193 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 194

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(120 , 8)) report "TEST FALLITO. Expected  120  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 194 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 195

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(106 , 8)) report "TEST FALLITO. Expected  106  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 195 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 196

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(76 , 8)) report "TEST FALLITO. Expected  76  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 196 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 197

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(4 , 8)) report "TEST FALLITO. Expected  4  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 197 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 198 interrotto

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		--interruzione dopo reset
		--tb_start <= '1';
		--wait for c_CLOCK_PERIOD;
		--wait until tb_done = '1';
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(20 , 8)) report "TEST FALLITO. Expected  20  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 198 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 199 asincrono

		wait for 600 ns;-----------------------attesa pi� lunga per colpire il componente durante uno stato diverso
		--wait for c_CLOCK_PERIOD;-------------test asincrono
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(107 , 8)) report "TEST FALLITO. Expected  107  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 199 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 200

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(58 , 8)) report "TEST FALLITO. Expected  58  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 200 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 201

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(129 , 8)) report "TEST FALLITO. Expected  129  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 201 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 202

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(116 , 8)) report "TEST FALLITO. Expected  116  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 202 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 203

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(129 , 8)) report "TEST FALLITO. Expected  129  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 203 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 204

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(212 , 8)) report "TEST FALLITO. Expected  212  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 204 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 205

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(31 , 8)) report "TEST FALLITO. Expected  31  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 205 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 206

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(200 , 8)) report "TEST FALLITO. Expected  200  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 206 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 207

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(117 , 8)) report "TEST FALLITO. Expected  117  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 207 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 208

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(34 , 8)) report "TEST FALLITO. Expected  34  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 208 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 209

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(28 , 8)) report "TEST FALLITO. Expected  28  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 209 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 210

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(98 , 8)) report "TEST FALLITO. Expected  98  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 210 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 211

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(6 , 8)) report "TEST FALLITO. Expected  6  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 211 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 212

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(60 , 8)) report "TEST FALLITO. Expected  60  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 212 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 213

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(161 , 8)) report "TEST FALLITO. Expected  161  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 213 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 214

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(22 , 8)) report "TEST FALLITO. Expected  22  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 214 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 215

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(216 , 8)) report "TEST FALLITO. Expected  216  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 215 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 216

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(28 , 8)) report "TEST FALLITO. Expected  28  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 216 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 217

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(49 , 8)) report "TEST FALLITO. Expected  49  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 217 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 218

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(209 , 8)) report "TEST FALLITO. Expected  209  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 218 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 219

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(27 , 8)) report "TEST FALLITO. Expected  27  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 219 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 220

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(43 , 8)) report "TEST FALLITO. Expected  43  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 220 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 221

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(178 , 8)) report "TEST FALLITO. Expected  178  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 221 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 222

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(74 , 8)) report "TEST FALLITO. Expected  74  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 222 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 223

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(106 , 8)) report "TEST FALLITO. Expected  106  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 223 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 224

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(25 , 8)) report "TEST FALLITO. Expected  25  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 224 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 225

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(118 , 8)) report "TEST FALLITO. Expected  118  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 225 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 226

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(127 , 8)) report "TEST FALLITO. Expected  127  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 226 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 227

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(33 , 8)) report "TEST FALLITO. Expected  33  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 227 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 228

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(0 , 8)) report "TEST FALLITO. Expected  0  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 228 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 229

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(132 , 8)) report "TEST FALLITO. Expected  132  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 229 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 230

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(20 , 8)) report "TEST FALLITO. Expected  20  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 230 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 231

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(7 , 8)) report "TEST FALLITO. Expected  7  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 231 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 232

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(5 , 8)) report "TEST FALLITO. Expected  5  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 232 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 233

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(145 , 8)) report "TEST FALLITO. Expected  145  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 233 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 234

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(43 , 8)) report "TEST FALLITO. Expected  43  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 234 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 235

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(177 , 8)) report "TEST FALLITO. Expected  177  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 235 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 236

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(145 , 8)) report "TEST FALLITO. Expected  145  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 236 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 237

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(89 , 8)) report "TEST FALLITO. Expected  89  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 237 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 238

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(216 , 8)) report "TEST FALLITO. Expected  216  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 238 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 239

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(248 , 8)) report "TEST FALLITO. Expected  248  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 239 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 240

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(95 , 8)) report "TEST FALLITO. Expected  95  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 240 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 241

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(13 , 8)) report "TEST FALLITO. Expected  13  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 241 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 242

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(79 , 8)) report "TEST FALLITO. Expected  79  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 242 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 243

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(12 , 8)) report "TEST FALLITO. Expected  12  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 243 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 244

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(64 , 8)) report "TEST FALLITO. Expected  64  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 244 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 245

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(48 , 8)) report "TEST FALLITO. Expected  48  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 245 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 246

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(98 , 8)) report "TEST FALLITO. Expected  98  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 246 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 247

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(52 , 8)) report "TEST FALLITO. Expected  52  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 247 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 248 interrotto

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		--interruzione
		--wait for c_CLOCK_PERIOD;
		--wait until tb_done = '1';
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(77 , 8)) report "TEST FALLITO. Expected  77  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 248 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 249 asincrono

		wait for 1000 ns;-------------------attesa diversa per colpire durante uno stato diverso
		--wait for c_CLOCK_PERIOD;----------test asincrono
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(52 , 8)) report "TEST FALLITO. Expected  52  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 249 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 250

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(59 , 8)) report "TEST FALLITO. Expected  59  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 250 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 251

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(77 , 8)) report "TEST FALLITO. Expected  77  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 251 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 252

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(112 , 8)) report "TEST FALLITO. Expected  112  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 252 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 253

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(52 , 8)) report "TEST FALLITO. Expected  52  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 253 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 254

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(72 , 8)) report "TEST FALLITO. Expected  72  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 254 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 255

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(42 , 8)) report "TEST FALLITO. Expected  42  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 255 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 256

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(80 , 8)) report "TEST FALLITO. Expected  80  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 256 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 257

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(23 , 8)) report "TEST FALLITO. Expected  23  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 257 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 258

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(120 , 8)) report "TEST FALLITO. Expected  120  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 258 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 259

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(3 , 8)) report "TEST FALLITO. Expected  3  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 259 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 260

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(129 , 8)) report "TEST FALLITO. Expected  129  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 260 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 261

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(74 , 8)) report "TEST FALLITO. Expected  74  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 261 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 262

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(122 , 8)) report "TEST FALLITO. Expected  122  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 262 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 263

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(117 , 8)) report "TEST FALLITO. Expected  117  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 263 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 264

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(193 , 8)) report "TEST FALLITO. Expected  193  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 264 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 265

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(244 , 8)) report "TEST FALLITO. Expected  244  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 265 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 266

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(241 , 8)) report "TEST FALLITO. Expected  241  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 266 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 267

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(98 , 8)) report "TEST FALLITO. Expected  98  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 267 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 268

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(97 , 8)) report "TEST FALLITO. Expected  97  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 268 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 269

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(72 , 8)) report "TEST FALLITO. Expected  72  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 269 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 270

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(57 , 8)) report "TEST FALLITO. Expected  57  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 270 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 271

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(109 , 8)) report "TEST FALLITO. Expected  109  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 271 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 272

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(212 , 8)) report "TEST FALLITO. Expected  212  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 272 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 273

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(105 , 8)) report "TEST FALLITO. Expected  105  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 273 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 274

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(26 , 8)) report "TEST FALLITO. Expected  26  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 274 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 275

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(4 , 8)) report "TEST FALLITO. Expected  4  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 275 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 276

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(244 , 8)) report "TEST FALLITO. Expected  244  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 276 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 277

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(125 , 8)) report "TEST FALLITO. Expected  125  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 277 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 278

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(118 , 8)) report "TEST FALLITO. Expected  118  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 278 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 279

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(111 , 8)) report "TEST FALLITO. Expected  111  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 279 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 280

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(74 , 8)) report "TEST FALLITO. Expected  74  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 280 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 281

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(148 , 8)) report "TEST FALLITO. Expected  148  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 281 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 282

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(47 , 8)) report "TEST FALLITO. Expected  47  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 282 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 283

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(59 , 8)) report "TEST FALLITO. Expected  59  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 283 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 284

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(152 , 8)) report "TEST FALLITO. Expected  152  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 284 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 285

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(83 , 8)) report "TEST FALLITO. Expected  83  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 285 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 286

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(152 , 8)) report "TEST FALLITO. Expected  152  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 286 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 287

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(42 , 8)) report "TEST FALLITO. Expected  42  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 287 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 288

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(41 , 8)) report "TEST FALLITO. Expected  41  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 288 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 289

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(178 , 8)) report "TEST FALLITO. Expected  178  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 289 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 290

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(67 , 8)) report "TEST FALLITO. Expected  67  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 290 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 291

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(108 , 8)) report "TEST FALLITO. Expected  108  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 291 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 292

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(226 , 8)) report "TEST FALLITO. Expected  226  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 292 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 293

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(34 , 8)) report "TEST FALLITO. Expected  34  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 293 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 294

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(92 , 8)) report "TEST FALLITO. Expected  92  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 294 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 295

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(75 , 8)) report "TEST FALLITO. Expected  75  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 295 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 296

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(123 , 8)) report "TEST FALLITO. Expected  123  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 296 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 297

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(83 , 8)) report "TEST FALLITO. Expected  83  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 297 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 298 interrotto. Saranno interrotti diversi test successivi per testare reset asincroni multipli

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		--interruzione
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(94 , 8)) report "TEST FALLITO. Expected  94  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 298 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 299 asincrono e interrotto

		wait for 300 ns;-----------------attesa non standard
		--wait for c_CLOCK_PERIOD;-------reset asincrono
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		--interruzione
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '1';
		--wait for c_CLOCK_PERIOD;
		--wait until tb_done = '1';
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(216 , 8)) report "TEST FALLITO. Expected  216  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 299 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 300 interrotto

		wait for 10 ns;------------------attesa non standard
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		--interruzione
		--wait for c_CLOCK_PERIOD;
		--wait until tb_done = '1';
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(56 , 8)) report "TEST FALLITO. Expected  56  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 300 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 301 asincrono e interrotto

		wait for 50 ns;--------------attesa non standard
		--wait for c_CLOCK_PERIOD;---reset asincrono
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		--interruzione 
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '1';
		--wait for c_CLOCK_PERIOD;
		--wait until tb_done = '1';
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(194 , 8)) report "TEST FALLITO. Expected  194  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 301 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 302 asincrono

		wait for 300 ns;------------attesa non standard
		--wait for c_CLOCK_PERIOD;--reset asincrono
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '1';----------start � alto da due reset fa
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(111 , 8)) report "TEST FALLITO. Expected  111  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 302 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 303

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(59 , 8)) report "TEST FALLITO. Expected  59  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 303 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 304

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(68 , 8)) report "TEST FALLITO. Expected  68  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 304 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 305

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(55 , 8)) report "TEST FALLITO. Expected  55  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 305 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 306

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(248 , 8)) report "TEST FALLITO. Expected  248  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 306 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 307

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(54 , 8)) report "TEST FALLITO. Expected  54  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 307 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 308

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(35 , 8)) report "TEST FALLITO. Expected  35  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 308 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 309

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(63 , 8)) report "TEST FALLITO. Expected  63  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 309 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 310

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(120 , 8)) report "TEST FALLITO. Expected  120  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 310 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 311

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(97 , 8)) report "TEST FALLITO. Expected  97  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 311 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 312

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(162 , 8)) report "TEST FALLITO. Expected  162  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 312 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 313

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(59 , 8)) report "TEST FALLITO. Expected  59  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 313 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 314

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(39 , 8)) report "TEST FALLITO. Expected  39  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 314 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 315

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(29 , 8)) report "TEST FALLITO. Expected  29  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 315 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 316

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(92 , 8)) report "TEST FALLITO. Expected  92  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 316 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 317

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(61 , 8)) report "TEST FALLITO. Expected  61  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 317 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 318

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(21 , 8)) report "TEST FALLITO. Expected  21  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 318 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 319

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(180 , 8)) report "TEST FALLITO. Expected  180  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 319 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 320

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(111 , 8)) report "TEST FALLITO. Expected  111  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 320 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 321

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(62 , 8)) report "TEST FALLITO. Expected  62  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 321 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 322

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(152 , 8)) report "TEST FALLITO. Expected  152  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 322 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 323

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(38 , 8)) report "TEST FALLITO. Expected  38  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 323 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 324

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(72 , 8)) report "TEST FALLITO. Expected  72  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 324 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 325

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(49 , 8)) report "TEST FALLITO. Expected  49  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 325 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 326

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(36 , 8)) report "TEST FALLITO. Expected  36  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 326 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 327

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(79 , 8)) report "TEST FALLITO. Expected  79  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 327 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 328

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(92 , 8)) report "TEST FALLITO. Expected  92  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 328 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 329

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(112 , 8)) report "TEST FALLITO. Expected  112  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 329 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 330

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(111 , 8)) report "TEST FALLITO. Expected  111  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 330 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 331

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(145 , 8)) report "TEST FALLITO. Expected  145  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 331 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 332

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(49 , 8)) report "TEST FALLITO. Expected  49  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 332 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 333

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(126 , 8)) report "TEST FALLITO. Expected  126  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 333 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 334

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(59 , 8)) report "TEST FALLITO. Expected  59  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 334 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 335

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(87 , 8)) report "TEST FALLITO. Expected  87  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 335 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 336

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(100 , 8)) report "TEST FALLITO. Expected  100  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 336 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 337

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(50 , 8)) report "TEST FALLITO. Expected  50  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 337 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 338

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(148 , 8)) report "TEST FALLITO. Expected  148  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 338 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 339

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(29 , 8)) report "TEST FALLITO. Expected  29  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 339 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 340

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(71 , 8)) report "TEST FALLITO. Expected  71  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 340 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 341

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(124 , 8)) report "TEST FALLITO. Expected  124  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 341 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 342

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(89 , 8)) report "TEST FALLITO. Expected  89  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 342 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 343

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(184 , 8)) report "TEST FALLITO. Expected  184  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 343 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 344

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(22 , 8)) report "TEST FALLITO. Expected  22  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 344 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 345

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(21 , 8)) report "TEST FALLITO. Expected  21  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 345 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 346

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(161 , 8)) report "TEST FALLITO. Expected  161  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 346 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 347

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(180 , 8)) report "TEST FALLITO. Expected  180  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 347 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 348 interrotto

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		--interruzione
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '1';
		--wait for c_CLOCK_PERIOD;
		--wait until tb_done = '1';
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(28 , 8)) report "TEST FALLITO. Expected  28  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 348 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 349 asincrono

		wait for 1 ns;--------------------attesa brevissima prima di nuovo reset
		--wait for c_CLOCK_PERIOD;--------reset asincrono
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(34 , 8)) report "TEST FALLITO. Expected  34  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 349 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 350

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(124 , 8)) report "TEST FALLITO. Expected  124  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 350 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 351

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(33 , 8)) report "TEST FALLITO. Expected  33  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 351 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 352

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(9 , 8)) report "TEST FALLITO. Expected  9  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 352 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 353

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(161 , 8)) report "TEST FALLITO. Expected  161  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 353 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 354

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(72 , 8)) report "TEST FALLITO. Expected  72  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 354 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 355

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(72 , 8)) report "TEST FALLITO. Expected  72  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 355 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 356

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(9 , 8)) report "TEST FALLITO. Expected  9  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 356 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 357

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(152 , 8)) report "TEST FALLITO. Expected  152  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 357 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 358

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(73 , 8)) report "TEST FALLITO. Expected  73  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 358 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 359

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(210 , 8)) report "TEST FALLITO. Expected  210  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 359 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 360

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(5 , 8)) report "TEST FALLITO. Expected  5  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 360 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 361

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(31 , 8)) report "TEST FALLITO. Expected  31  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 361 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 362

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(116 , 8)) report "TEST FALLITO. Expected  116  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 362 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 363

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(110 , 8)) report "TEST FALLITO. Expected  110  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 363 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 364

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(27 , 8)) report "TEST FALLITO. Expected  27  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 364 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 365

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(125 , 8)) report "TEST FALLITO. Expected  125  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 365 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 366

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(132 , 8)) report "TEST FALLITO. Expected  132  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 366 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 367

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(241 , 8)) report "TEST FALLITO. Expected  241  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 367 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 368

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(145 , 8)) report "TEST FALLITO. Expected  145  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 368 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 369

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(83 , 8)) report "TEST FALLITO. Expected  83  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 369 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 370

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(10 , 8)) report "TEST FALLITO. Expected  10  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 370 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 371

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(31 , 8)) report "TEST FALLITO. Expected  31  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 371 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 372

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(164 , 8)) report "TEST FALLITO. Expected  164  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 372 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 373

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(82 , 8)) report "TEST FALLITO. Expected  82  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 373 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 374

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(61 , 8)) report "TEST FALLITO. Expected  61  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 374 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 375

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(36 , 8)) report "TEST FALLITO. Expected  36  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 375 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 376

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(8 , 8)) report "TEST FALLITO. Expected  8  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 376 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 377

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(161 , 8)) report "TEST FALLITO. Expected  161  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 377 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 378

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(110 , 8)) report "TEST FALLITO. Expected  110  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 378 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 379

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(108 , 8)) report "TEST FALLITO. Expected  108  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 379 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 380

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(29 , 8)) report "TEST FALLITO. Expected  29  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 380 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 381

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(113 , 8)) report "TEST FALLITO. Expected  113  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 381 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 382

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(145 , 8)) report "TEST FALLITO. Expected  145  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 382 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 383

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(177 , 8)) report "TEST FALLITO. Expected  177  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 383 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 384

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(146 , 8)) report "TEST FALLITO. Expected  146  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 384 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 385

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(35 , 8)) report "TEST FALLITO. Expected  35  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 385 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 386

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(26 , 8)) report "TEST FALLITO. Expected  26  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 386 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 387

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(46 , 8)) report "TEST FALLITO. Expected  46  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 387 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 388

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(127 , 8)) report "TEST FALLITO. Expected  127  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 388 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 389

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(95 , 8)) report "TEST FALLITO. Expected  95  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 389 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 390

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(161 , 8)) report "TEST FALLITO. Expected  161  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 390 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 391

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(40 , 8)) report "TEST FALLITO. Expected  40  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 391 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 392

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(86 , 8)) report "TEST FALLITO. Expected  86  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 392 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 393

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(13 , 8)) report "TEST FALLITO. Expected  13  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 393 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 394

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(225 , 8)) report "TEST FALLITO. Expected  225  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 394 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 395

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(8 , 8)) report "TEST FALLITO. Expected  8  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 395 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 396

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(25 , 8)) report "TEST FALLITO. Expected  25  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 396 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 397

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(120 , 8)) report "TEST FALLITO. Expected  120  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 397 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 398 interrotto

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		--interruzione
		--wait for c_CLOCK_PERIOD;
		--wait until tb_done = '1';
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(244 , 8)) report "TEST FALLITO. Expected  244  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 398 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 399 asincrono

		wait for 5000 ns;--------------------attesa molto lunga dopo start
		--wait for c_CLOCK_PERIOD;-----------reset asincrono
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		--tb_start <= '1';-------------------alto dal test precedente
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(90 , 8)) report "TEST FALLITO. Expected  90  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 399 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 400

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(29 , 8)) report "TEST FALLITO. Expected  29  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 400 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 401

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(226 , 8)) report "TEST FALLITO. Expected  226  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 401 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 402

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(130 , 8)) report "TEST FALLITO. Expected  130  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 402 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 403

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(209 , 8)) report "TEST FALLITO. Expected  209  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 403 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 404

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(107 , 8)) report "TEST FALLITO. Expected  107  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 404 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 405

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(32 , 8)) report "TEST FALLITO. Expected  32  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 405 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 406

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(85 , 8)) report "TEST FALLITO. Expected  85  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 406 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 407

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(118 , 8)) report "TEST FALLITO. Expected  118  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 407 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 408

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(168 , 8)) report "TEST FALLITO. Expected  168  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 408 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 409

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(129 , 8)) report "TEST FALLITO. Expected  129  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 409 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 410

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(178 , 8)) report "TEST FALLITO. Expected  178  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 410 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 411

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(61 , 8)) report "TEST FALLITO. Expected  61  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 411 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 412

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(85 , 8)) report "TEST FALLITO. Expected  85  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 412 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 413

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(78 , 8)) report "TEST FALLITO. Expected  78  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 413 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 414

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(60 , 8)) report "TEST FALLITO. Expected  60  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 414 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 415

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(4 , 8)) report "TEST FALLITO. Expected  4  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 415 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 416

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(136 , 8)) report "TEST FALLITO. Expected  136  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 416 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 417

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(121 , 8)) report "TEST FALLITO. Expected  121  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 417 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 418

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(57 , 8)) report "TEST FALLITO. Expected  57  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 418 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 419

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(17 , 8)) report "TEST FALLITO. Expected  17  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 419 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 420

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(27 , 8)) report "TEST FALLITO. Expected  27  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 420 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 421

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(0 , 8)) report "TEST FALLITO. Expected  0  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 421 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 422

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(51 , 8)) report "TEST FALLITO. Expected  51  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 422 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 423

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(117 , 8)) report "TEST FALLITO. Expected  117  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 423 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 424

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(210 , 8)) report "TEST FALLITO. Expected  210  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 424 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 425

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(42 , 8)) report "TEST FALLITO. Expected  42  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 425 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 426

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(96 , 8)) report "TEST FALLITO. Expected  96  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 426 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 427

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(76 , 8)) report "TEST FALLITO. Expected  76  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 427 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 428

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(46 , 8)) report "TEST FALLITO. Expected  46  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 428 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 429

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(117 , 8)) report "TEST FALLITO. Expected  117  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 429 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 430

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(232 , 8)) report "TEST FALLITO. Expected  232  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 430 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 431

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(77 , 8)) report "TEST FALLITO. Expected  77  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 431 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 432

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(12 , 8)) report "TEST FALLITO. Expected  12  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 432 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 433

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(76 , 8)) report "TEST FALLITO. Expected  76  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 433 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 434

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(117 , 8)) report "TEST FALLITO. Expected  117  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 434 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 435

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(162 , 8)) report "TEST FALLITO. Expected  162  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 435 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 436

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(118 , 8)) report "TEST FALLITO. Expected  118  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 436 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 437

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(45 , 8)) report "TEST FALLITO. Expected  45  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 437 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 438

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(228 , 8)) report "TEST FALLITO. Expected  228  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 438 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 439

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(56 , 8)) report "TEST FALLITO. Expected  56  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 439 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 440

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(125 , 8)) report "TEST FALLITO. Expected  125  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 440 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 441

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(107 , 8)) report "TEST FALLITO. Expected  107  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 441 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 442

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(12 , 8)) report "TEST FALLITO. Expected  12  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 442 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 443

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(59 , 8)) report "TEST FALLITO. Expected  59  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 443 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 444

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(24 , 8)) report "TEST FALLITO. Expected  24  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 444 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 445

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(42 , 8)) report "TEST FALLITO. Expected  42  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 445 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 446

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(45 , 8)) report "TEST FALLITO. Expected  45  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 446 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 447

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(50 , 8)) report "TEST FALLITO. Expected  50  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 447 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 448 interrotto

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';-----------------start alzato prima di reset
		tb_rst <= '0';
		
		--interruzione
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '1';
		--wait for c_CLOCK_PERIOD;
		--wait until tb_done = '1';
		--wait for c_CLOCK_PERIOD;
		--tb_start <= '0';
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(212 , 8)) report "TEST FALLITO. Expected  212  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 448 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 449 asincrono

		wait for 10 ns;--------------------------attesa breve
		--wait for c_CLOCK_PERIOD;---------------reset asincrono
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		--tb_start <= '1';-----------------------alto da prima
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(79 , 8)) report "TEST FALLITO. Expected  79  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 449 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 450

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(110 , 8)) report "TEST FALLITO. Expected  110  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 450 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 451

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(78 , 8)) report "TEST FALLITO. Expected  78  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 451 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 452

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(216 , 8)) report "TEST FALLITO. Expected  216  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 452 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 453

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(226 , 8)) report "TEST FALLITO. Expected  226  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 453 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 454

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(62 , 8)) report "TEST FALLITO. Expected  62  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 454 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 455

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(18 , 8)) report "TEST FALLITO. Expected  18  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 455 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 456

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(42 , 8)) report "TEST FALLITO. Expected  42  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 456 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 457

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(85 , 8)) report "TEST FALLITO. Expected  85  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 457 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 458

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(45 , 8)) report "TEST FALLITO. Expected  45  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 458 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 459

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(111 , 8)) report "TEST FALLITO. Expected  111  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 459 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 460

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(37 , 8)) report "TEST FALLITO. Expected  37  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 460 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 461

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(67 , 8)) report "TEST FALLITO. Expected  67  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 461 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 462

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(19 , 8)) report "TEST FALLITO. Expected  19  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 462 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 463

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(59 , 8)) report "TEST FALLITO. Expected  59  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 463 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 464

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(164 , 8)) report "TEST FALLITO. Expected  164  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 464 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 465

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(94 , 8)) report "TEST FALLITO. Expected  94  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 465 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 466

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(30 , 8)) report "TEST FALLITO. Expected  30  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 466 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 467

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(39 , 8)) report "TEST FALLITO. Expected  39  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 467 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 468

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(5 , 8)) report "TEST FALLITO. Expected  5  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 468 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 469

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(65 , 8)) report "TEST FALLITO. Expected  65  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 469 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 470

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(232 , 8)) report "TEST FALLITO. Expected  232  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 470 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 471

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(95 , 8)) report "TEST FALLITO. Expected  95  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 471 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 472

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(105 , 8)) report "TEST FALLITO. Expected  105  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 472 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 473

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(40 , 8)) report "TEST FALLITO. Expected  40  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 473 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 474

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(93 , 8)) report "TEST FALLITO. Expected  93  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 474 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 475

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(61 , 8)) report "TEST FALLITO. Expected  61  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 475 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 476

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(184 , 8)) report "TEST FALLITO. Expected  184  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 476 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 477

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(28 , 8)) report "TEST FALLITO. Expected  28  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 477 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 478

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(148 , 8)) report "TEST FALLITO. Expected  148  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 478 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 479

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(7 , 8)) report "TEST FALLITO. Expected  7  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 479 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 480

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(216 , 8)) report "TEST FALLITO. Expected  216  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 480 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 481

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(161 , 8)) report "TEST FALLITO. Expected  161  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 481 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 482

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(125 , 8)) report "TEST FALLITO. Expected  125  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 482 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 483

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(225 , 8)) report "TEST FALLITO. Expected  225  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 483 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 484

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(8 , 8)) report "TEST FALLITO. Expected  8  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 484 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 485

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(61 , 8)) report "TEST FALLITO. Expected  61  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 485 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 486

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(106 , 8)) report "TEST FALLITO. Expected  106  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 486 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 487

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(93 , 8)) report "TEST FALLITO. Expected  93  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 487 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 488

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(248 , 8)) report "TEST FALLITO. Expected  248  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 488 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 489

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(57 , 8)) report "TEST FALLITO. Expected  57  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 489 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 490

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(193 , 8)) report "TEST FALLITO. Expected  193  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 490 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 491

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(26 , 8)) report "TEST FALLITO. Expected  26  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 491 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 492

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(130 , 8)) report "TEST FALLITO. Expected  130  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 492 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 493

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(180 , 8)) report "TEST FALLITO. Expected  180  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 493 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 494

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(52 , 8)) report "TEST FALLITO. Expected  52  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 494 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 495

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(126 , 8)) report "TEST FALLITO. Expected  126  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 495 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 496

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(36 , 8)) report "TEST FALLITO. Expected  36  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 496 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 497

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(52 , 8)) report "TEST FALLITO. Expected  52  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 497 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 498 interrotto

		wait for 100 ns;
		wait for c_CLOCK_PERIOD;
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		--interruzione
		--wait until tb_done = '0';
		--wait for 100 ns;

		--assert RAM(9) = std_logic_vector(to_unsigned(196 , 8)) report "TEST FALLITO. Expected  196  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		--report "TEST 498 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		-- test numero 499

		wait for 10 ns;
		--wait for c_CLOCK_PERIOD;------------------reset asincrono
		tb_rst <= '1';
		wait for c_CLOCK_PERIOD;
		tb_rst <= '0';
		wait for c_CLOCK_PERIOD;
		tb_start <= '1';
		wait for c_CLOCK_PERIOD;
		wait until tb_done = '1';
		wait for c_CLOCK_PERIOD;
		tb_start <= '0';
		wait until tb_done = '0';
		wait for 100 ns;

		assert RAM(9) = std_logic_vector(to_unsigned(106 , 8)) report "TEST FALLITO. Expected  106  found " & integer'image(to_integer(unsigned(RAM(9))))  severity failure;

		report "TEST 499 PASSATO sol: " & integer'image(to_integer(unsigned(RAM(9))));


		assert false report "TUTTO OK"  severity failure;
	end process test;
end projecttb;
